/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 18:59:13 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1478065269 */

module registerNbits__0_18(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module registerNbits__0_21(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module datapath(b_mantissa, a_mantissa, o_mantissa);
   input [23:0]b_mantissa;
   input [23:0]a_mantissa;
   output [47:0]o_mantissa;

   HA_X1 i_0 (.A(n_1494), .B(n_1785), .CO(n_1), .S(n_0));
   FA_X1 i_1 (.A(n_1471), .B(n_1493), .CI(n_1515), .CO(n_3), .S(n_2));
   HA_X1 i_2 (.A(n_1535), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_3 (.A(n_1448), .B(n_1470), .CI(n_1492), .CO(n_7), .S(n_6));
   FA_X1 i_4 (.A(n_1514), .B(n_1534), .CI(n_5), .CO(n_9), .S(n_8));
   HA_X1 i_5 (.A(n_3), .B(n_8), .CO(n_11), .S(n_10));
   FA_X1 i_6 (.A(n_1425), .B(n_1447), .CI(n_1469), .CO(n_13), .S(n_12));
   FA_X1 i_7 (.A(n_1491), .B(n_1513), .CI(n_1533), .CO(n_15), .S(n_14));
   FA_X1 i_8 (.A(n_7), .B(n_9), .CI(n_14), .CO(n_17), .S(n_16));
   HA_X1 i_9 (.A(n_12), .B(n_11), .CO(n_19), .S(n_18));
   FA_X1 i_10 (.A(n_1402), .B(n_1424), .CI(n_1446), .CO(n_21), .S(n_20));
   FA_X1 i_11 (.A(n_1468), .B(n_1490), .CI(n_1512), .CO(n_23), .S(n_22));
   FA_X1 i_12 (.A(n_1532), .B(n_15), .CI(n_13), .CO(n_25), .S(n_24));
   FA_X1 i_13 (.A(n_22), .B(n_20), .CI(n_24), .CO(n_27), .S(n_26));
   HA_X1 i_14 (.A(n_19), .B(n_17), .CO(n_29), .S(n_28));
   FA_X1 i_15 (.A(n_1379), .B(n_1401), .CI(n_1423), .CO(n_31), .S(n_30));
   FA_X1 i_16 (.A(n_1445), .B(n_1467), .CI(n_1489), .CO(n_33), .S(n_32));
   FA_X1 i_17 (.A(n_1511), .B(n_1531), .CI(n_23), .CO(n_35), .S(n_34));
   FA_X1 i_18 (.A(n_21), .B(n_25), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_19 (.A(n_32), .B(n_30), .CI(n_29), .CO(n_39), .S(n_38));
   HA_X1 i_20 (.A(n_36), .B(n_27), .CO(n_41), .S(n_40));
   FA_X1 i_21 (.A(n_1356), .B(n_1378), .CI(n_1400), .CO(n_43), .S(n_42));
   FA_X1 i_22 (.A(n_1422), .B(n_1444), .CI(n_1466), .CO(n_45), .S(n_44));
   FA_X1 i_23 (.A(n_1488), .B(n_1510), .CI(n_1530), .CO(n_47), .S(n_46));
   FA_X1 i_24 (.A(n_33), .B(n_31), .CI(n_35), .CO(n_49), .S(n_48));
   FA_X1 i_25 (.A(n_46), .B(n_44), .CI(n_42), .CO(n_51), .S(n_50));
   FA_X1 i_26 (.A(n_48), .B(n_37), .CI(n_41), .CO(n_53), .S(n_52));
   HA_X1 i_27 (.A(n_39), .B(n_50), .CO(n_55), .S(n_54));
   FA_X1 i_28 (.A(n_1333), .B(n_1355), .CI(n_1377), .CO(n_57), .S(n_56));
   FA_X1 i_29 (.A(n_1399), .B(n_1421), .CI(n_1443), .CO(n_59), .S(n_58));
   FA_X1 i_30 (.A(n_1465), .B(n_1487), .CI(n_1509), .CO(n_61), .S(n_60));
   FA_X1 i_31 (.A(n_1529), .B(n_47), .CI(n_45), .CO(n_63), .S(n_62));
   FA_X1 i_32 (.A(n_43), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_33 (.A(n_56), .B(n_49), .CI(n_62), .CO(n_67), .S(n_66));
   FA_X1 i_34 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_35 (.A(n_55), .B(n_53), .CO(n_71), .S(n_70));
   FA_X1 i_36 (.A(n_1310), .B(n_1332), .CI(n_1354), .CO(n_73), .S(n_72));
   FA_X1 i_37 (.A(n_1376), .B(n_1398), .CI(n_1420), .CO(n_75), .S(n_74));
   FA_X1 i_38 (.A(n_1442), .B(n_1464), .CI(n_1486), .CO(n_77), .S(n_76));
   FA_X1 i_39 (.A(n_1508), .B(n_1528), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_40 (.A(n_59), .B(n_57), .CI(n_63), .CO(n_81), .S(n_80));
   FA_X1 i_41 (.A(n_78), .B(n_76), .CI(n_74), .CO(n_83), .S(n_82));
   FA_X1 i_42 (.A(n_72), .B(n_80), .CI(n_65), .CO(n_85), .S(n_84));
   FA_X1 i_43 (.A(n_67), .B(n_82), .CI(n_84), .CO(n_87), .S(n_86));
   HA_X1 i_44 (.A(n_71), .B(n_69), .CO(n_89), .S(n_88));
   FA_X1 i_45 (.A(n_1287), .B(n_1309), .CI(n_1331), .CO(n_91), .S(n_90));
   FA_X1 i_46 (.A(n_1353), .B(n_1375), .CI(n_1397), .CO(n_93), .S(n_92));
   FA_X1 i_47 (.A(n_1419), .B(n_1441), .CI(n_1463), .CO(n_95), .S(n_94));
   FA_X1 i_48 (.A(n_1485), .B(n_1507), .CI(n_1527), .CO(n_97), .S(n_96));
   FA_X1 i_49 (.A(n_77), .B(n_75), .CI(n_73), .CO(n_99), .S(n_98));
   FA_X1 i_50 (.A(n_79), .B(n_96), .CI(n_94), .CO(n_101), .S(n_100));
   FA_X1 i_51 (.A(n_92), .B(n_90), .CI(n_81), .CO(n_103), .S(n_102));
   FA_X1 i_52 (.A(n_98), .B(n_83), .CI(n_85), .CO(n_105), .S(n_104));
   FA_X1 i_53 (.A(n_102), .B(n_100), .CI(n_104), .CO(n_107), .S(n_106));
   HA_X1 i_54 (.A(n_89), .B(n_87), .CO(n_109), .S(n_108));
   FA_X1 i_55 (.A(n_1264), .B(n_1286), .CI(n_1308), .CO(n_111), .S(n_110));
   FA_X1 i_56 (.A(n_1330), .B(n_1352), .CI(n_1374), .CO(n_113), .S(n_112));
   FA_X1 i_57 (.A(n_1396), .B(n_1418), .CI(n_1440), .CO(n_115), .S(n_114));
   FA_X1 i_58 (.A(n_1462), .B(n_1484), .CI(n_1506), .CO(n_117), .S(n_116));
   FA_X1 i_59 (.A(n_1526), .B(n_97), .CI(n_95), .CO(n_119), .S(n_118));
   FA_X1 i_60 (.A(n_93), .B(n_91), .CI(n_99), .CO(n_121), .S(n_120));
   FA_X1 i_61 (.A(n_116), .B(n_114), .CI(n_112), .CO(n_123), .S(n_122));
   FA_X1 i_62 (.A(n_110), .B(n_120), .CI(n_118), .CO(n_125), .S(n_124));
   FA_X1 i_63 (.A(n_101), .B(n_103), .CI(n_122), .CO(n_127), .S(n_126));
   FA_X1 i_64 (.A(n_105), .B(n_124), .CI(n_126), .CO(n_129), .S(n_128));
   HA_X1 i_65 (.A(n_107), .B(n_109), .CO(n_131), .S(n_130));
   FA_X1 i_66 (.A(n_1241), .B(n_1263), .CI(n_1285), .CO(n_133), .S(n_132));
   FA_X1 i_67 (.A(n_1307), .B(n_1329), .CI(n_1351), .CO(n_135), .S(n_134));
   FA_X1 i_68 (.A(n_1373), .B(n_1395), .CI(n_1417), .CO(n_137), .S(n_136));
   FA_X1 i_69 (.A(n_1439), .B(n_1461), .CI(n_1483), .CO(n_139), .S(n_138));
   FA_X1 i_70 (.A(n_1505), .B(n_1525), .CI(n_117), .CO(n_141), .S(n_140));
   FA_X1 i_71 (.A(n_115), .B(n_113), .CI(n_111), .CO(n_143), .S(n_142));
   FA_X1 i_72 (.A(n_119), .B(n_140), .CI(n_138), .CO(n_145), .S(n_144));
   FA_X1 i_73 (.A(n_136), .B(n_134), .CI(n_132), .CO(n_147), .S(n_146));
   FA_X1 i_74 (.A(n_121), .B(n_142), .CI(n_123), .CO(n_149), .S(n_148));
   FA_X1 i_75 (.A(n_125), .B(n_146), .CI(n_144), .CO(n_151), .S(n_150));
   FA_X1 i_76 (.A(n_148), .B(n_127), .CI(n_129), .CO(n_153), .S(n_152));
   HA_X1 i_77 (.A(n_150), .B(n_131), .CO(n_155), .S(n_154));
   FA_X1 i_78 (.A(n_1218), .B(n_1240), .CI(n_1262), .CO(n_157), .S(n_156));
   FA_X1 i_79 (.A(n_1284), .B(n_1306), .CI(n_1328), .CO(n_159), .S(n_158));
   FA_X1 i_80 (.A(n_1350), .B(n_1372), .CI(n_1394), .CO(n_161), .S(n_160));
   FA_X1 i_81 (.A(n_1416), .B(n_1438), .CI(n_1460), .CO(n_163), .S(n_162));
   FA_X1 i_82 (.A(n_1482), .B(n_1504), .CI(n_1524), .CO(n_165), .S(n_164));
   FA_X1 i_83 (.A(n_139), .B(n_137), .CI(n_135), .CO(n_167), .S(n_166));
   FA_X1 i_84 (.A(n_133), .B(n_143), .CI(n_141), .CO(n_169), .S(n_168));
   FA_X1 i_85 (.A(n_164), .B(n_162), .CI(n_160), .CO(n_171), .S(n_170));
   FA_X1 i_86 (.A(n_158), .B(n_156), .CI(n_166), .CO(n_173), .S(n_172));
   FA_X1 i_87 (.A(n_147), .B(n_145), .CI(n_168), .CO(n_175), .S(n_174));
   FA_X1 i_88 (.A(n_149), .B(n_172), .CI(n_170), .CO(n_177), .S(n_176));
   FA_X1 i_89 (.A(n_174), .B(n_151), .CI(n_176), .CO(n_179), .S(n_178));
   HA_X1 i_90 (.A(n_153), .B(n_155), .CO(n_181), .S(n_180));
   FA_X1 i_91 (.A(n_1195), .B(n_1217), .CI(n_1239), .CO(n_183), .S(n_182));
   FA_X1 i_92 (.A(n_1261), .B(n_1283), .CI(n_1305), .CO(n_185), .S(n_184));
   FA_X1 i_93 (.A(n_1327), .B(n_1349), .CI(n_1371), .CO(n_187), .S(n_186));
   FA_X1 i_94 (.A(n_1393), .B(n_1415), .CI(n_1437), .CO(n_189), .S(n_188));
   FA_X1 i_95 (.A(n_1459), .B(n_1481), .CI(n_1503), .CO(n_191), .S(n_190));
   FA_X1 i_96 (.A(n_1523), .B(n_165), .CI(n_163), .CO(n_193), .S(n_192));
   FA_X1 i_97 (.A(n_161), .B(n_159), .CI(n_157), .CO(n_195), .S(n_194));
   FA_X1 i_98 (.A(n_167), .B(n_190), .CI(n_188), .CO(n_197), .S(n_196));
   FA_X1 i_99 (.A(n_186), .B(n_184), .CI(n_182), .CO(n_199), .S(n_198));
   FA_X1 i_100 (.A(n_169), .B(n_194), .CI(n_192), .CO(n_201), .S(n_200));
   FA_X1 i_101 (.A(n_171), .B(n_173), .CI(n_198), .CO(n_203), .S(n_202));
   FA_X1 i_102 (.A(n_196), .B(n_175), .CI(n_200), .CO(n_205), .S(n_204));
   FA_X1 i_103 (.A(n_177), .B(n_202), .CI(n_204), .CO(n_207), .S(n_206));
   HA_X1 i_104 (.A(n_179), .B(n_181), .CO(n_209), .S(n_208));
   FA_X1 i_105 (.A(n_1172), .B(n_1194), .CI(n_1216), .CO(n_211), .S(n_210));
   FA_X1 i_106 (.A(n_1238), .B(n_1260), .CI(n_1282), .CO(n_213), .S(n_212));
   FA_X1 i_107 (.A(n_1304), .B(n_1326), .CI(n_1348), .CO(n_215), .S(n_214));
   FA_X1 i_108 (.A(n_1370), .B(n_1392), .CI(n_1414), .CO(n_217), .S(n_216));
   FA_X1 i_109 (.A(n_1436), .B(n_1458), .CI(n_1480), .CO(n_219), .S(n_218));
   FA_X1 i_110 (.A(n_1502), .B(n_1522), .CI(n_191), .CO(n_221), .S(n_220));
   FA_X1 i_111 (.A(n_189), .B(n_187), .CI(n_185), .CO(n_223), .S(n_222));
   FA_X1 i_112 (.A(n_183), .B(n_195), .CI(n_193), .CO(n_225), .S(n_224));
   FA_X1 i_113 (.A(n_220), .B(n_218), .CI(n_216), .CO(n_227), .S(n_226));
   FA_X1 i_114 (.A(n_214), .B(n_212), .CI(n_210), .CO(n_229), .S(n_228));
   FA_X1 i_115 (.A(n_222), .B(n_199), .CI(n_197), .CO(n_231), .S(n_230));
   FA_X1 i_116 (.A(n_224), .B(n_201), .CI(n_228), .CO(n_233), .S(n_232));
   FA_X1 i_117 (.A(n_226), .B(n_230), .CI(n_203), .CO(n_235), .S(n_234));
   FA_X1 i_118 (.A(n_232), .B(n_205), .CI(n_234), .CO(n_237), .S(n_236));
   HA_X1 i_119 (.A(n_207), .B(n_209), .CO(n_239), .S(n_238));
   FA_X1 i_120 (.A(n_1149), .B(n_1171), .CI(n_1193), .CO(n_241), .S(n_240));
   FA_X1 i_121 (.A(n_1215), .B(n_1237), .CI(n_1259), .CO(n_243), .S(n_242));
   FA_X1 i_122 (.A(n_1281), .B(n_1303), .CI(n_1325), .CO(n_245), .S(n_244));
   FA_X1 i_123 (.A(n_1347), .B(n_1369), .CI(n_1391), .CO(n_247), .S(n_246));
   FA_X1 i_124 (.A(n_1413), .B(n_1435), .CI(n_1457), .CO(n_249), .S(n_248));
   FA_X1 i_125 (.A(n_1479), .B(n_1501), .CI(n_1521), .CO(n_251), .S(n_250));
   FA_X1 i_126 (.A(n_219), .B(n_217), .CI(n_215), .CO(n_253), .S(n_252));
   FA_X1 i_127 (.A(n_213), .B(n_211), .CI(n_223), .CO(n_255), .S(n_254));
   FA_X1 i_128 (.A(n_221), .B(n_250), .CI(n_248), .CO(n_257), .S(n_256));
   FA_X1 i_129 (.A(n_246), .B(n_244), .CI(n_242), .CO(n_259), .S(n_258));
   FA_X1 i_130 (.A(n_240), .B(n_225), .CI(n_254), .CO(n_261), .S(n_260));
   FA_X1 i_131 (.A(n_252), .B(n_229), .CI(n_227), .CO(n_263), .S(n_262));
   FA_X1 i_132 (.A(n_231), .B(n_258), .CI(n_256), .CO(n_265), .S(n_264));
   FA_X1 i_133 (.A(n_260), .B(n_262), .CI(n_233), .CO(n_267), .S(n_266));
   FA_X1 i_134 (.A(n_235), .B(n_264), .CI(n_266), .CO(n_269), .S(n_268));
   HA_X1 i_135 (.A(n_237), .B(n_239), .CO(n_271), .S(n_270));
   FA_X1 i_136 (.A(n_1126), .B(n_1148), .CI(n_1170), .CO(n_273), .S(n_272));
   FA_X1 i_137 (.A(n_1192), .B(n_1214), .CI(n_1236), .CO(n_275), .S(n_274));
   FA_X1 i_138 (.A(n_1258), .B(n_1280), .CI(n_1302), .CO(n_277), .S(n_276));
   FA_X1 i_139 (.A(n_1324), .B(n_1346), .CI(n_1368), .CO(n_279), .S(n_278));
   FA_X1 i_140 (.A(n_1390), .B(n_1412), .CI(n_1434), .CO(n_281), .S(n_280));
   FA_X1 i_141 (.A(n_1456), .B(n_1478), .CI(n_1500), .CO(n_283), .S(n_282));
   FA_X1 i_142 (.A(n_1520), .B(n_251), .CI(n_249), .CO(n_285), .S(n_284));
   FA_X1 i_143 (.A(n_247), .B(n_245), .CI(n_243), .CO(n_287), .S(n_286));
   FA_X1 i_144 (.A(n_241), .B(n_253), .CI(n_282), .CO(n_289), .S(n_288));
   FA_X1 i_145 (.A(n_280), .B(n_278), .CI(n_276), .CO(n_291), .S(n_290));
   FA_X1 i_146 (.A(n_274), .B(n_272), .CI(n_255), .CO(n_293), .S(n_292));
   FA_X1 i_147 (.A(n_286), .B(n_284), .CI(n_259), .CO(n_295), .S(n_294));
   FA_X1 i_148 (.A(n_257), .B(n_288), .CI(n_263), .CO(n_297), .S(n_296));
   FA_X1 i_149 (.A(n_261), .B(n_292), .CI(n_290), .CO(n_299), .S(n_298));
   FA_X1 i_150 (.A(n_294), .B(n_265), .CI(n_296), .CO(n_301), .S(n_300));
   FA_X1 i_151 (.A(n_267), .B(n_298), .CI(n_300), .CO(n_303), .S(n_302));
   HA_X1 i_152 (.A(n_269), .B(n_302), .CO(n_305), .S(n_304));
   FA_X1 i_153 (.A(n_1103), .B(n_1125), .CI(n_1147), .CO(n_307), .S(n_306));
   FA_X1 i_154 (.A(n_1169), .B(n_1191), .CI(n_1213), .CO(n_309), .S(n_308));
   FA_X1 i_155 (.A(n_1235), .B(n_1257), .CI(n_1279), .CO(n_311), .S(n_310));
   FA_X1 i_156 (.A(n_1301), .B(n_1323), .CI(n_1345), .CO(n_313), .S(n_312));
   FA_X1 i_157 (.A(n_1367), .B(n_1389), .CI(n_1411), .CO(n_315), .S(n_314));
   FA_X1 i_158 (.A(n_1433), .B(n_1455), .CI(n_1477), .CO(n_317), .S(n_316));
   FA_X1 i_159 (.A(n_1499), .B(n_1519), .CI(n_283), .CO(n_319), .S(n_318));
   FA_X1 i_160 (.A(n_281), .B(n_279), .CI(n_277), .CO(n_321), .S(n_320));
   FA_X1 i_161 (.A(n_275), .B(n_273), .CI(n_287), .CO(n_323), .S(n_322));
   FA_X1 i_162 (.A(n_285), .B(n_318), .CI(n_316), .CO(n_325), .S(n_324));
   FA_X1 i_163 (.A(n_314), .B(n_312), .CI(n_310), .CO(n_327), .S(n_326));
   FA_X1 i_164 (.A(n_308), .B(n_306), .CI(n_322), .CO(n_329), .S(n_328));
   FA_X1 i_165 (.A(n_320), .B(n_291), .CI(n_289), .CO(n_331), .S(n_330));
   FA_X1 i_166 (.A(n_293), .B(n_295), .CI(n_328), .CO(n_333), .S(n_332));
   FA_X1 i_167 (.A(n_326), .B(n_324), .CI(n_297), .CO(n_335), .S(n_334));
   FA_X1 i_168 (.A(n_330), .B(n_299), .CI(n_332), .CO(n_337), .S(n_336));
   FA_X1 i_169 (.A(n_334), .B(n_301), .CI(n_336), .CO(n_339), .S(n_338));
   HA_X1 i_170 (.A(n_303), .B(n_338), .CO(n_341), .S(n_340));
   FA_X1 i_171 (.A(n_1080), .B(n_1102), .CI(n_1124), .CO(n_343), .S(n_342));
   FA_X1 i_172 (.A(n_1146), .B(n_1168), .CI(n_1190), .CO(n_345), .S(n_344));
   FA_X1 i_173 (.A(n_1212), .B(n_1234), .CI(n_1256), .CO(n_347), .S(n_346));
   FA_X1 i_174 (.A(n_1278), .B(n_1300), .CI(n_1322), .CO(n_349), .S(n_348));
   FA_X1 i_175 (.A(n_1344), .B(n_1366), .CI(n_1388), .CO(n_351), .S(n_350));
   FA_X1 i_176 (.A(n_1410), .B(n_1432), .CI(n_1454), .CO(n_353), .S(n_352));
   FA_X1 i_177 (.A(n_1476), .B(n_1498), .CI(n_1518), .CO(n_355), .S(n_354));
   FA_X1 i_178 (.A(n_317), .B(n_315), .CI(n_313), .CO(n_357), .S(n_356));
   FA_X1 i_179 (.A(n_311), .B(n_309), .CI(n_307), .CO(n_359), .S(n_358));
   FA_X1 i_180 (.A(n_321), .B(n_319), .CI(n_354), .CO(n_361), .S(n_360));
   FA_X1 i_181 (.A(n_352), .B(n_350), .CI(n_348), .CO(n_363), .S(n_362));
   FA_X1 i_182 (.A(n_346), .B(n_344), .CI(n_342), .CO(n_365), .S(n_364));
   FA_X1 i_183 (.A(n_323), .B(n_358), .CI(n_356), .CO(n_367), .S(n_366));
   FA_X1 i_184 (.A(n_327), .B(n_325), .CI(n_360), .CO(n_369), .S(n_368));
   FA_X1 i_185 (.A(n_331), .B(n_329), .CI(n_364), .CO(n_371), .S(n_370));
   FA_X1 i_186 (.A(n_362), .B(n_368), .CI(n_366), .CO(n_373), .S(n_372));
   FA_X1 i_187 (.A(n_333), .B(n_335), .CI(n_370), .CO(n_375), .S(n_374));
   FA_X1 i_188 (.A(n_337), .B(n_372), .CI(n_374), .CO(n_377), .S(n_376));
   HA_X1 i_189 (.A(n_339), .B(n_341), .CO(n_379), .S(n_378));
   FA_X1 i_190 (.A(n_1057), .B(n_1079), .CI(n_1101), .CO(n_381), .S(n_380));
   FA_X1 i_191 (.A(n_1123), .B(n_1145), .CI(n_1167), .CO(n_383), .S(n_382));
   FA_X1 i_192 (.A(n_1189), .B(n_1211), .CI(n_1233), .CO(n_385), .S(n_384));
   FA_X1 i_193 (.A(n_1255), .B(n_1277), .CI(n_1299), .CO(n_387), .S(n_386));
   FA_X1 i_194 (.A(n_1321), .B(n_1343), .CI(n_1365), .CO(n_389), .S(n_388));
   FA_X1 i_195 (.A(n_1387), .B(n_1409), .CI(n_1431), .CO(n_391), .S(n_390));
   FA_X1 i_196 (.A(n_1453), .B(n_1475), .CI(n_1497), .CO(n_393), .S(n_392));
   FA_X1 i_197 (.A(n_1517), .B(n_355), .CI(n_353), .CO(n_395), .S(n_394));
   FA_X1 i_198 (.A(n_351), .B(n_349), .CI(n_347), .CO(n_397), .S(n_396));
   FA_X1 i_199 (.A(n_345), .B(n_343), .CI(n_359), .CO(n_399), .S(n_398));
   FA_X1 i_200 (.A(n_357), .B(n_392), .CI(n_390), .CO(n_401), .S(n_400));
   FA_X1 i_201 (.A(n_388), .B(n_386), .CI(n_384), .CO(n_403), .S(n_402));
   FA_X1 i_202 (.A(n_382), .B(n_380), .CI(n_398), .CO(n_405), .S(n_404));
   FA_X1 i_203 (.A(n_396), .B(n_394), .CI(n_365), .CO(n_407), .S(n_406));
   FA_X1 i_204 (.A(n_363), .B(n_361), .CI(n_367), .CO(n_409), .S(n_408));
   FA_X1 i_205 (.A(n_404), .B(n_402), .CI(n_400), .CO(n_411), .S(n_410));
   FA_X1 i_206 (.A(n_369), .B(n_408), .CI(n_406), .CO(n_413), .S(n_412));
   FA_X1 i_207 (.A(n_371), .B(n_373), .CI(n_410), .CO(n_415), .S(n_414));
   FA_X1 i_208 (.A(n_375), .B(n_412), .CI(n_414), .CO(n_417), .S(n_416));
   HA_X1 i_209 (.A(n_377), .B(n_416), .CO(n_419), .S(n_418));
   FA_X1 i_210 (.A(n_1034), .B(n_1056), .CI(n_1078), .CO(n_421), .S(n_420));
   FA_X1 i_211 (.A(n_1100), .B(n_1122), .CI(n_1144), .CO(n_423), .S(n_422));
   FA_X1 i_212 (.A(n_1166), .B(n_1188), .CI(n_1210), .CO(n_425), .S(n_424));
   FA_X1 i_213 (.A(n_1232), .B(n_1254), .CI(n_1276), .CO(n_427), .S(n_426));
   FA_X1 i_214 (.A(n_1298), .B(n_1320), .CI(n_1342), .CO(n_429), .S(n_428));
   FA_X1 i_215 (.A(n_1364), .B(n_1386), .CI(n_1408), .CO(n_431), .S(n_430));
   FA_X1 i_216 (.A(n_1430), .B(n_1452), .CI(n_1474), .CO(n_433), .S(n_432));
   FA_X1 i_217 (.A(n_1496), .B(n_1516), .CI(n_393), .CO(n_435), .S(n_434));
   FA_X1 i_218 (.A(n_391), .B(n_389), .CI(n_387), .CO(n_437), .S(n_436));
   FA_X1 i_219 (.A(n_385), .B(n_383), .CI(n_381), .CO(n_439), .S(n_438));
   FA_X1 i_220 (.A(n_397), .B(n_395), .CI(n_434), .CO(n_441), .S(n_440));
   FA_X1 i_221 (.A(n_432), .B(n_430), .CI(n_428), .CO(n_443), .S(n_442));
   FA_X1 i_222 (.A(n_426), .B(n_424), .CI(n_422), .CO(n_445), .S(n_444));
   FA_X1 i_223 (.A(n_420), .B(n_399), .CI(n_438), .CO(n_447), .S(n_446));
   FA_X1 i_224 (.A(n_436), .B(n_403), .CI(n_401), .CO(n_449), .S(n_448));
   FA_X1 i_225 (.A(n_440), .B(n_407), .CI(n_405), .CO(n_451), .S(n_450));
   FA_X1 i_226 (.A(n_444), .B(n_442), .CI(n_446), .CO(n_453), .S(n_452));
   FA_X1 i_227 (.A(n_409), .B(n_448), .CI(n_411), .CO(n_455), .S(n_454));
   FA_X1 i_228 (.A(n_450), .B(n_413), .CI(n_452), .CO(n_457), .S(n_456));
   FA_X1 i_229 (.A(n_454), .B(n_415), .CI(n_456), .CO(n_459), .S(n_458));
   HA_X1 i_230 (.A(n_417), .B(n_458), .CO(n_461), .S(n_460));
   FA_X1 i_231 (.A(a_mantissa[0]), .B(n_1033), .CI(n_1055), .CO(n_463), .S(n_462));
   FA_X1 i_232 (.A(n_1077), .B(n_1099), .CI(n_1121), .CO(n_465), .S(n_464));
   FA_X1 i_233 (.A(n_1143), .B(n_1165), .CI(n_1187), .CO(n_467), .S(n_466));
   FA_X1 i_234 (.A(n_1209), .B(n_1231), .CI(n_1253), .CO(n_469), .S(n_468));
   FA_X1 i_235 (.A(n_1275), .B(n_1297), .CI(n_1319), .CO(n_471), .S(n_470));
   FA_X1 i_236 (.A(n_1341), .B(n_1363), .CI(n_1385), .CO(n_473), .S(n_472));
   FA_X1 i_237 (.A(n_1407), .B(n_1429), .CI(n_1451), .CO(n_475), .S(n_474));
   FA_X1 i_238 (.A(n_1473), .B(n_1495), .CI(b_mantissa[0]), .CO(n_477), .S(n_476));
   FA_X1 i_239 (.A(n_433), .B(n_431), .CI(n_429), .CO(n_479), .S(n_478));
   FA_X1 i_240 (.A(n_427), .B(n_425), .CI(n_423), .CO(n_481), .S(n_480));
   FA_X1 i_241 (.A(n_421), .B(n_439), .CI(n_437), .CO(n_483), .S(n_482));
   FA_X1 i_242 (.A(n_435), .B(n_476), .CI(n_474), .CO(n_485), .S(n_484));
   FA_X1 i_243 (.A(n_472), .B(n_470), .CI(n_468), .CO(n_487), .S(n_486));
   FA_X1 i_244 (.A(n_466), .B(n_464), .CI(n_462), .CO(n_489), .S(n_488));
   FA_X1 i_245 (.A(n_480), .B(n_478), .CI(n_445), .CO(n_491), .S(n_490));
   FA_X1 i_246 (.A(n_443), .B(n_441), .CI(n_482), .CO(n_493), .S(n_492));
   FA_X1 i_247 (.A(n_449), .B(n_447), .CI(n_488), .CO(n_495), .S(n_494));
   FA_X1 i_248 (.A(n_486), .B(n_484), .CI(n_451), .CO(n_497), .S(n_496));
   FA_X1 i_249 (.A(n_492), .B(n_490), .CI(n_453), .CO(n_499), .S(n_498));
   FA_X1 i_250 (.A(n_494), .B(n_455), .CI(n_496), .CO(n_501), .S(n_500));
   FA_X1 i_251 (.A(n_498), .B(n_457), .CI(n_500), .CO(n_503), .S(n_502));
   HA_X1 i_252 (.A(n_459), .B(n_502), .CO(n_505), .S(n_504));
   FA_X1 i_253 (.A(a_mantissa[1]), .B(n_1032), .CI(n_1054), .CO(n_507), .S(n_506));
   FA_X1 i_254 (.A(n_1076), .B(n_1098), .CI(n_1120), .CO(n_509), .S(n_508));
   FA_X1 i_255 (.A(n_1142), .B(n_1164), .CI(n_1186), .CO(n_511), .S(n_510));
   FA_X1 i_256 (.A(n_1208), .B(n_1230), .CI(n_1252), .CO(n_513), .S(n_512));
   FA_X1 i_257 (.A(n_1274), .B(n_1296), .CI(n_1318), .CO(n_515), .S(n_514));
   FA_X1 i_258 (.A(n_1340), .B(n_1362), .CI(n_1384), .CO(n_517), .S(n_516));
   FA_X1 i_259 (.A(n_1406), .B(n_1428), .CI(n_1450), .CO(n_519), .S(n_518));
   FA_X1 i_260 (.A(n_1472), .B(b_mantissa[1]), .CI(n_477), .CO(n_521), .S(n_520));
   FA_X1 i_261 (.A(n_475), .B(n_473), .CI(n_471), .CO(n_523), .S(n_522));
   FA_X1 i_262 (.A(n_469), .B(n_467), .CI(n_465), .CO(n_525), .S(n_524));
   FA_X1 i_263 (.A(n_463), .B(n_481), .CI(n_479), .CO(n_527), .S(n_526));
   FA_X1 i_264 (.A(n_520), .B(n_518), .CI(n_516), .CO(n_529), .S(n_528));
   FA_X1 i_265 (.A(n_514), .B(n_512), .CI(n_510), .CO(n_531), .S(n_530));
   FA_X1 i_266 (.A(n_508), .B(n_506), .CI(n_483), .CO(n_533), .S(n_532));
   FA_X1 i_267 (.A(n_524), .B(n_522), .CI(n_489), .CO(n_535), .S(n_534));
   FA_X1 i_268 (.A(n_487), .B(n_485), .CI(n_526), .CO(n_537), .S(n_536));
   FA_X1 i_269 (.A(n_491), .B(n_532), .CI(n_530), .CO(n_539), .S(n_538));
   FA_X1 i_270 (.A(n_528), .B(n_493), .CI(n_536), .CO(n_541), .S(n_540));
   FA_X1 i_271 (.A(n_534), .B(n_495), .CI(n_497), .CO(n_543), .S(n_542));
   FA_X1 i_272 (.A(n_499), .B(n_538), .CI(n_540), .CO(n_545), .S(n_544));
   FA_X1 i_273 (.A(n_542), .B(n_501), .CI(n_544), .CO(n_547), .S(n_546));
   HA_X1 i_274 (.A(n_503), .B(n_546), .CO(n_549), .S(n_548));
   FA_X1 i_275 (.A(a_mantissa[2]), .B(n_1031), .CI(n_1053), .CO(n_551), .S(n_550));
   FA_X1 i_276 (.A(n_1075), .B(n_1097), .CI(n_1119), .CO(n_553), .S(n_552));
   FA_X1 i_277 (.A(n_1141), .B(n_1163), .CI(n_1185), .CO(n_555), .S(n_554));
   FA_X1 i_278 (.A(n_1207), .B(n_1229), .CI(n_1251), .CO(n_557), .S(n_556));
   FA_X1 i_279 (.A(n_1273), .B(n_1295), .CI(n_1317), .CO(n_559), .S(n_558));
   FA_X1 i_280 (.A(n_1339), .B(n_1361), .CI(n_1383), .CO(n_561), .S(n_560));
   FA_X1 i_281 (.A(n_1405), .B(n_1427), .CI(n_1449), .CO(n_563), .S(n_562));
   FA_X1 i_282 (.A(b_mantissa[2]), .B(n_519), .CI(n_517), .CO(n_565), .S(n_564));
   FA_X1 i_283 (.A(n_515), .B(n_513), .CI(n_511), .CO(n_567), .S(n_566));
   FA_X1 i_284 (.A(n_509), .B(n_507), .CI(n_525), .CO(n_569), .S(n_568));
   FA_X1 i_285 (.A(n_523), .B(n_521), .CI(n_562), .CO(n_571), .S(n_570));
   FA_X1 i_286 (.A(n_560), .B(n_558), .CI(n_556), .CO(n_573), .S(n_572));
   FA_X1 i_287 (.A(n_554), .B(n_552), .CI(n_550), .CO(n_575), .S(n_574));
   FA_X1 i_288 (.A(n_527), .B(n_568), .CI(n_566), .CO(n_577), .S(n_576));
   FA_X1 i_289 (.A(n_564), .B(n_531), .CI(n_529), .CO(n_579), .S(n_578));
   FA_X1 i_290 (.A(n_533), .B(n_570), .CI(n_535), .CO(n_581), .S(n_580));
   FA_X1 i_291 (.A(n_574), .B(n_572), .CI(n_537), .CO(n_583), .S(n_582));
   FA_X1 i_292 (.A(n_578), .B(n_576), .CI(n_539), .CO(n_585), .S(n_584));
   FA_X1 i_293 (.A(n_580), .B(n_541), .CI(n_543), .CO(n_587), .S(n_586));
   FA_X1 i_294 (.A(n_582), .B(n_584), .CI(n_545), .CO(n_589), .S(n_588));
   FA_X1 i_295 (.A(n_586), .B(n_588), .CI(n_547), .CO(n_591), .S(n_590));
   FA_X1 i_296 (.A(a_mantissa[3]), .B(n_1030), .CI(n_1052), .CO(n_593), .S(n_592));
   FA_X1 i_297 (.A(n_1074), .B(n_1096), .CI(n_1118), .CO(n_595), .S(n_594));
   FA_X1 i_298 (.A(n_1140), .B(n_1162), .CI(n_1184), .CO(n_597), .S(n_596));
   FA_X1 i_299 (.A(n_1206), .B(n_1228), .CI(n_1250), .CO(n_599), .S(n_598));
   FA_X1 i_300 (.A(n_1272), .B(n_1294), .CI(n_1316), .CO(n_601), .S(n_600));
   FA_X1 i_301 (.A(n_1338), .B(n_1360), .CI(n_1382), .CO(n_603), .S(n_602));
   FA_X1 i_302 (.A(n_1404), .B(n_1426), .CI(b_mantissa[3]), .CO(n_605), .S(n_604));
   FA_X1 i_303 (.A(n_563), .B(n_561), .CI(n_559), .CO(n_607), .S(n_606));
   FA_X1 i_304 (.A(n_557), .B(n_555), .CI(n_553), .CO(n_609), .S(n_608));
   FA_X1 i_305 (.A(n_551), .B(n_567), .CI(n_565), .CO(n_611), .S(n_610));
   FA_X1 i_306 (.A(n_604), .B(n_602), .CI(n_600), .CO(n_613), .S(n_612));
   FA_X1 i_307 (.A(n_598), .B(n_596), .CI(n_594), .CO(n_615), .S(n_614));
   FA_X1 i_308 (.A(n_592), .B(n_569), .CI(n_608), .CO(n_617), .S(n_616));
   FA_X1 i_309 (.A(n_606), .B(n_575), .CI(n_573), .CO(n_619), .S(n_618));
   FA_X1 i_310 (.A(n_571), .B(n_610), .CI(n_579), .CO(n_621), .S(n_620));
   FA_X1 i_311 (.A(n_577), .B(n_614), .CI(n_612), .CO(n_623), .S(n_622));
   FA_X1 i_312 (.A(n_616), .B(n_581), .CI(n_618), .CO(n_625), .S(n_624));
   FA_X1 i_313 (.A(n_583), .B(n_620), .CI(n_585), .CO(n_627), .S(n_626));
   FA_X1 i_314 (.A(n_622), .B(n_624), .CI(n_587), .CO(n_629), .S(n_628));
   FA_X1 i_315 (.A(n_626), .B(n_589), .CI(n_628), .CO(n_631), .S(n_630));
   FA_X1 i_316 (.A(a_mantissa[4]), .B(n_1029), .CI(n_1051), .CO(n_633), .S(n_632));
   FA_X1 i_317 (.A(n_1073), .B(n_1095), .CI(n_1117), .CO(n_635), .S(n_634));
   FA_X1 i_318 (.A(n_1139), .B(n_1161), .CI(n_1183), .CO(n_637), .S(n_636));
   FA_X1 i_319 (.A(n_1205), .B(n_1227), .CI(n_1249), .CO(n_639), .S(n_638));
   FA_X1 i_320 (.A(n_1271), .B(n_1293), .CI(n_1315), .CO(n_641), .S(n_640));
   FA_X1 i_321 (.A(n_1337), .B(n_1359), .CI(n_1381), .CO(n_643), .S(n_642));
   FA_X1 i_322 (.A(n_1403), .B(b_mantissa[4]), .CI(n_605), .CO(n_645), .S(n_644));
   FA_X1 i_323 (.A(n_603), .B(n_601), .CI(n_599), .CO(n_647), .S(n_646));
   FA_X1 i_324 (.A(n_597), .B(n_595), .CI(n_593), .CO(n_649), .S(n_648));
   FA_X1 i_325 (.A(n_609), .B(n_607), .CI(n_644), .CO(n_651), .S(n_650));
   FA_X1 i_326 (.A(n_642), .B(n_640), .CI(n_638), .CO(n_653), .S(n_652));
   FA_X1 i_327 (.A(n_636), .B(n_634), .CI(n_632), .CO(n_655), .S(n_654));
   FA_X1 i_328 (.A(n_611), .B(n_648), .CI(n_646), .CO(n_657), .S(n_656));
   FA_X1 i_329 (.A(n_615), .B(n_613), .CI(n_650), .CO(n_659), .S(n_658));
   FA_X1 i_330 (.A(n_619), .B(n_617), .CI(n_654), .CO(n_661), .S(n_660));
   FA_X1 i_331 (.A(n_652), .B(n_621), .CI(n_658), .CO(n_663), .S(n_662));
   FA_X1 i_332 (.A(n_656), .B(n_623), .CI(n_660), .CO(n_665), .S(n_664));
   FA_X1 i_333 (.A(n_625), .B(n_662), .CI(n_627), .CO(n_667), .S(n_666));
   FA_X1 i_334 (.A(n_664), .B(n_629), .CI(n_666), .CO(n_669), .S(n_668));
   FA_X1 i_335 (.A(a_mantissa[5]), .B(n_1028), .CI(n_1050), .CO(n_671), .S(n_670));
   FA_X1 i_336 (.A(n_1072), .B(n_1094), .CI(n_1116), .CO(n_673), .S(n_672));
   FA_X1 i_337 (.A(n_1138), .B(n_1160), .CI(n_1182), .CO(n_675), .S(n_674));
   FA_X1 i_338 (.A(n_1204), .B(n_1226), .CI(n_1248), .CO(n_677), .S(n_676));
   FA_X1 i_339 (.A(n_1270), .B(n_1292), .CI(n_1314), .CO(n_679), .S(n_678));
   FA_X1 i_340 (.A(n_1336), .B(n_1358), .CI(n_1380), .CO(n_681), .S(n_680));
   FA_X1 i_341 (.A(b_mantissa[5]), .B(n_643), .CI(n_641), .CO(n_683), .S(n_682));
   FA_X1 i_342 (.A(n_639), .B(n_637), .CI(n_635), .CO(n_685), .S(n_684));
   FA_X1 i_343 (.A(n_633), .B(n_649), .CI(n_647), .CO(n_687), .S(n_686));
   FA_X1 i_344 (.A(n_645), .B(n_680), .CI(n_678), .CO(n_689), .S(n_688));
   FA_X1 i_345 (.A(n_676), .B(n_674), .CI(n_672), .CO(n_691), .S(n_690));
   FA_X1 i_346 (.A(n_670), .B(n_684), .CI(n_682), .CO(n_693), .S(n_692));
   FA_X1 i_347 (.A(n_655), .B(n_653), .CI(n_651), .CO(n_695), .S(n_694));
   FA_X1 i_348 (.A(n_686), .B(n_657), .CI(n_690), .CO(n_697), .S(n_696));
   FA_X1 i_349 (.A(n_688), .B(n_659), .CI(n_694), .CO(n_699), .S(n_698));
   FA_X1 i_350 (.A(n_692), .B(n_661), .CI(n_696), .CO(n_701), .S(n_700));
   FA_X1 i_351 (.A(n_663), .B(n_698), .CI(n_665), .CO(n_703), .S(n_702));
   FA_X1 i_352 (.A(n_700), .B(n_667), .CI(n_702), .CO(n_705), .S(n_704));
   FA_X1 i_353 (.A(a_mantissa[6]), .B(n_1027), .CI(n_1049), .CO(n_707), .S(n_706));
   FA_X1 i_354 (.A(n_1071), .B(n_1093), .CI(n_1115), .CO(n_709), .S(n_708));
   FA_X1 i_355 (.A(n_1137), .B(n_1159), .CI(n_1181), .CO(n_711), .S(n_710));
   FA_X1 i_356 (.A(n_1203), .B(n_1225), .CI(n_1247), .CO(n_713), .S(n_712));
   FA_X1 i_357 (.A(n_1269), .B(n_1291), .CI(n_1313), .CO(n_715), .S(n_714));
   FA_X1 i_358 (.A(n_1335), .B(n_1357), .CI(b_mantissa[6]), .CO(n_717), .S(n_716));
   FA_X1 i_359 (.A(n_681), .B(n_679), .CI(n_677), .CO(n_719), .S(n_718));
   FA_X1 i_360 (.A(n_675), .B(n_673), .CI(n_671), .CO(n_721), .S(n_720));
   FA_X1 i_361 (.A(n_685), .B(n_683), .CI(n_716), .CO(n_723), .S(n_722));
   FA_X1 i_362 (.A(n_714), .B(n_712), .CI(n_710), .CO(n_725), .S(n_724));
   FA_X1 i_363 (.A(n_708), .B(n_706), .CI(n_687), .CO(n_727), .S(n_726));
   FA_X1 i_364 (.A(n_720), .B(n_718), .CI(n_691), .CO(n_729), .S(n_728));
   FA_X1 i_365 (.A(n_689), .B(n_722), .CI(n_695), .CO(n_731), .S(n_730));
   FA_X1 i_366 (.A(n_693), .B(n_726), .CI(n_724), .CO(n_733), .S(n_732));
   FA_X1 i_367 (.A(n_728), .B(n_697), .CI(n_730), .CO(n_735), .S(n_734));
   FA_X1 i_368 (.A(n_699), .B(n_732), .CI(n_701), .CO(n_737), .S(n_736));
   FA_X1 i_369 (.A(n_734), .B(n_703), .CI(n_736), .CO(n_739), .S(n_738));
   FA_X1 i_370 (.A(a_mantissa[7]), .B(n_1026), .CI(n_1048), .CO(n_741), .S(n_740));
   FA_X1 i_371 (.A(n_1070), .B(n_1092), .CI(n_1114), .CO(n_743), .S(n_742));
   FA_X1 i_372 (.A(n_1136), .B(n_1158), .CI(n_1180), .CO(n_745), .S(n_744));
   FA_X1 i_373 (.A(n_1202), .B(n_1224), .CI(n_1246), .CO(n_747), .S(n_746));
   FA_X1 i_374 (.A(n_1268), .B(n_1290), .CI(n_1312), .CO(n_749), .S(n_748));
   FA_X1 i_375 (.A(n_1334), .B(b_mantissa[7]), .CI(n_717), .CO(n_751), .S(n_750));
   FA_X1 i_376 (.A(n_715), .B(n_713), .CI(n_711), .CO(n_753), .S(n_752));
   FA_X1 i_377 (.A(n_709), .B(n_707), .CI(n_721), .CO(n_755), .S(n_754));
   FA_X1 i_378 (.A(n_719), .B(n_750), .CI(n_748), .CO(n_757), .S(n_756));
   FA_X1 i_379 (.A(n_746), .B(n_744), .CI(n_742), .CO(n_759), .S(n_758));
   FA_X1 i_380 (.A(n_740), .B(n_754), .CI(n_752), .CO(n_761), .S(n_760));
   FA_X1 i_381 (.A(n_725), .B(n_723), .CI(n_727), .CO(n_763), .S(n_762));
   FA_X1 i_382 (.A(n_729), .B(n_758), .CI(n_756), .CO(n_765), .S(n_764));
   FA_X1 i_383 (.A(n_731), .B(n_762), .CI(n_760), .CO(n_767), .S(n_766));
   FA_X1 i_384 (.A(n_733), .B(n_764), .CI(n_735), .CO(n_769), .S(n_768));
   FA_X1 i_385 (.A(n_766), .B(n_737), .CI(n_768), .CO(n_771), .S(n_770));
   FA_X1 i_386 (.A(a_mantissa[8]), .B(n_1025), .CI(n_1047), .CO(n_773), .S(n_772));
   FA_X1 i_387 (.A(n_1069), .B(n_1091), .CI(n_1113), .CO(n_775), .S(n_774));
   FA_X1 i_388 (.A(n_1135), .B(n_1157), .CI(n_1179), .CO(n_777), .S(n_776));
   FA_X1 i_389 (.A(n_1201), .B(n_1223), .CI(n_1245), .CO(n_779), .S(n_778));
   FA_X1 i_390 (.A(n_1267), .B(n_1289), .CI(n_1311), .CO(n_781), .S(n_780));
   FA_X1 i_391 (.A(b_mantissa[8]), .B(n_749), .CI(n_747), .CO(n_783), .S(n_782));
   FA_X1 i_392 (.A(n_745), .B(n_743), .CI(n_741), .CO(n_785), .S(n_784));
   FA_X1 i_393 (.A(n_753), .B(n_751), .CI(n_780), .CO(n_787), .S(n_786));
   FA_X1 i_394 (.A(n_778), .B(n_776), .CI(n_774), .CO(n_789), .S(n_788));
   FA_X1 i_395 (.A(n_772), .B(n_755), .CI(n_784), .CO(n_791), .S(n_790));
   FA_X1 i_396 (.A(n_782), .B(n_759), .CI(n_757), .CO(n_793), .S(n_792));
   FA_X1 i_397 (.A(n_786), .B(n_761), .CI(n_763), .CO(n_795), .S(n_794));
   FA_X1 i_398 (.A(n_788), .B(n_790), .CI(n_792), .CO(n_797), .S(n_796));
   FA_X1 i_399 (.A(n_765), .B(n_794), .CI(n_767), .CO(n_799), .S(n_798));
   FA_X1 i_400 (.A(n_796), .B(n_769), .CI(n_798), .CO(n_801), .S(n_800));
   FA_X1 i_401 (.A(a_mantissa[9]), .B(n_1024), .CI(n_1046), .CO(n_803), .S(n_802));
   FA_X1 i_402 (.A(n_1068), .B(n_1090), .CI(n_1112), .CO(n_805), .S(n_804));
   FA_X1 i_403 (.A(n_1134), .B(n_1156), .CI(n_1178), .CO(n_807), .S(n_806));
   FA_X1 i_404 (.A(n_1200), .B(n_1222), .CI(n_1244), .CO(n_809), .S(n_808));
   FA_X1 i_405 (.A(n_1266), .B(n_1288), .CI(b_mantissa[9]), .CO(n_811), .S(n_810));
   FA_X1 i_406 (.A(n_781), .B(n_779), .CI(n_777), .CO(n_813), .S(n_812));
   FA_X1 i_407 (.A(n_775), .B(n_773), .CI(n_785), .CO(n_815), .S(n_814));
   FA_X1 i_408 (.A(n_783), .B(n_810), .CI(n_808), .CO(n_817), .S(n_816));
   FA_X1 i_409 (.A(n_806), .B(n_804), .CI(n_802), .CO(n_819), .S(n_818));
   FA_X1 i_410 (.A(n_814), .B(n_812), .CI(n_789), .CO(n_821), .S(n_820));
   FA_X1 i_411 (.A(n_787), .B(n_793), .CI(n_791), .CO(n_823), .S(n_822));
   FA_X1 i_412 (.A(n_818), .B(n_816), .CI(n_795), .CO(n_825), .S(n_824));
   FA_X1 i_413 (.A(n_820), .B(n_822), .CI(n_797), .CO(n_827), .S(n_826));
   FA_X1 i_414 (.A(n_824), .B(n_799), .CI(n_826), .CO(n_829), .S(n_828));
   FA_X1 i_415 (.A(a_mantissa[10]), .B(n_1023), .CI(n_1045), .CO(n_831), 
      .S(n_830));
   FA_X1 i_416 (.A(n_1067), .B(n_1089), .CI(n_1111), .CO(n_833), .S(n_832));
   FA_X1 i_417 (.A(n_1133), .B(n_1155), .CI(n_1177), .CO(n_835), .S(n_834));
   FA_X1 i_418 (.A(n_1199), .B(n_1221), .CI(n_1243), .CO(n_837), .S(n_836));
   FA_X1 i_419 (.A(n_1265), .B(b_mantissa[10]), .CI(n_811), .CO(n_839), .S(n_838));
   FA_X1 i_420 (.A(n_809), .B(n_807), .CI(n_805), .CO(n_841), .S(n_840));
   FA_X1 i_421 (.A(n_803), .B(n_813), .CI(n_838), .CO(n_843), .S(n_842));
   FA_X1 i_422 (.A(n_836), .B(n_834), .CI(n_832), .CO(n_845), .S(n_844));
   FA_X1 i_423 (.A(n_830), .B(n_815), .CI(n_840), .CO(n_847), .S(n_846));
   FA_X1 i_424 (.A(n_819), .B(n_817), .CI(n_842), .CO(n_849), .S(n_848));
   FA_X1 i_425 (.A(n_821), .B(n_844), .CI(n_846), .CO(n_851), .S(n_850));
   FA_X1 i_426 (.A(n_823), .B(n_848), .CI(n_825), .CO(n_853), .S(n_852));
   FA_X1 i_427 (.A(n_850), .B(n_827), .CI(n_852), .CO(n_855), .S(n_854));
   FA_X1 i_428 (.A(a_mantissa[11]), .B(n_1022), .CI(n_1044), .CO(n_857), 
      .S(n_856));
   FA_X1 i_429 (.A(n_1066), .B(n_1088), .CI(n_1110), .CO(n_859), .S(n_858));
   FA_X1 i_430 (.A(n_1132), .B(n_1154), .CI(n_1176), .CO(n_861), .S(n_860));
   FA_X1 i_431 (.A(n_1198), .B(n_1220), .CI(n_1242), .CO(n_863), .S(n_862));
   FA_X1 i_432 (.A(b_mantissa[11]), .B(n_837), .CI(n_835), .CO(n_865), .S(n_864));
   FA_X1 i_433 (.A(n_833), .B(n_831), .CI(n_841), .CO(n_867), .S(n_866));
   FA_X1 i_434 (.A(n_839), .B(n_862), .CI(n_860), .CO(n_869), .S(n_868));
   FA_X1 i_435 (.A(n_858), .B(n_856), .CI(n_866), .CO(n_871), .S(n_870));
   FA_X1 i_436 (.A(n_864), .B(n_845), .CI(n_843), .CO(n_873), .S(n_872));
   FA_X1 i_437 (.A(n_847), .B(n_870), .CI(n_868), .CO(n_875), .S(n_874));
   FA_X1 i_438 (.A(n_849), .B(n_872), .CI(n_851), .CO(n_877), .S(n_876));
   FA_X1 i_439 (.A(n_853), .B(n_874), .CI(n_876), .CO(n_879), .S(n_878));
   FA_X1 i_440 (.A(a_mantissa[12]), .B(n_1021), .CI(n_1043), .CO(n_881), 
      .S(n_880));
   FA_X1 i_441 (.A(n_1065), .B(n_1087), .CI(n_1109), .CO(n_883), .S(n_882));
   FA_X1 i_442 (.A(n_1131), .B(n_1153), .CI(n_1175), .CO(n_885), .S(n_884));
   FA_X1 i_443 (.A(n_1197), .B(n_1219), .CI(b_mantissa[12]), .CO(n_887), 
      .S(n_886));
   FA_X1 i_444 (.A(n_863), .B(n_861), .CI(n_859), .CO(n_889), .S(n_888));
   FA_X1 i_445 (.A(n_857), .B(n_865), .CI(n_886), .CO(n_891), .S(n_890));
   FA_X1 i_446 (.A(n_884), .B(n_882), .CI(n_880), .CO(n_893), .S(n_892));
   FA_X1 i_447 (.A(n_867), .B(n_888), .CI(n_869), .CO(n_895), .S(n_894));
   FA_X1 i_448 (.A(n_890), .B(n_873), .CI(n_871), .CO(n_897), .S(n_896));
   FA_X1 i_449 (.A(n_892), .B(n_894), .CI(n_875), .CO(n_899), .S(n_898));
   FA_X1 i_450 (.A(n_896), .B(n_877), .CI(n_898), .CO(n_901), .S(n_900));
   FA_X1 i_451 (.A(a_mantissa[13]), .B(n_1020), .CI(n_1042), .CO(n_903), 
      .S(n_902));
   FA_X1 i_452 (.A(n_1064), .B(n_1086), .CI(n_1108), .CO(n_905), .S(n_904));
   FA_X1 i_453 (.A(n_1130), .B(n_1152), .CI(n_1174), .CO(n_907), .S(n_906));
   FA_X1 i_454 (.A(n_1196), .B(b_mantissa[13]), .CI(n_887), .CO(n_909), .S(n_908));
   FA_X1 i_455 (.A(n_885), .B(n_883), .CI(n_881), .CO(n_911), .S(n_910));
   FA_X1 i_456 (.A(n_889), .B(n_908), .CI(n_906), .CO(n_913), .S(n_912));
   FA_X1 i_457 (.A(n_904), .B(n_902), .CI(n_910), .CO(n_915), .S(n_914));
   FA_X1 i_458 (.A(n_893), .B(n_891), .CI(n_895), .CO(n_917), .S(n_916));
   FA_X1 i_459 (.A(n_914), .B(n_912), .CI(n_897), .CO(n_919), .S(n_918));
   FA_X1 i_460 (.A(n_916), .B(n_899), .CI(n_918), .CO(n_921), .S(n_920));
   FA_X1 i_461 (.A(a_mantissa[14]), .B(n_1019), .CI(n_1041), .CO(n_923), 
      .S(n_922));
   FA_X1 i_462 (.A(n_1063), .B(n_1085), .CI(n_1107), .CO(n_925), .S(n_924));
   FA_X1 i_463 (.A(n_1129), .B(n_1151), .CI(n_1173), .CO(n_927), .S(n_926));
   FA_X1 i_464 (.A(b_mantissa[14]), .B(n_907), .CI(n_905), .CO(n_929), .S(n_928));
   FA_X1 i_465 (.A(n_903), .B(n_911), .CI(n_909), .CO(n_931), .S(n_930));
   FA_X1 i_466 (.A(n_926), .B(n_924), .CI(n_922), .CO(n_933), .S(n_932));
   FA_X1 i_467 (.A(n_928), .B(n_913), .CI(n_930), .CO(n_935), .S(n_934));
   FA_X1 i_468 (.A(n_915), .B(n_932), .CI(n_917), .CO(n_937), .S(n_936));
   FA_X1 i_469 (.A(n_934), .B(n_919), .CI(n_936), .CO(n_939), .S(n_938));
   FA_X1 i_470 (.A(a_mantissa[15]), .B(n_1018), .CI(n_1040), .CO(n_941), 
      .S(n_940));
   FA_X1 i_471 (.A(n_1062), .B(n_1084), .CI(n_1106), .CO(n_943), .S(n_942));
   FA_X1 i_472 (.A(n_1128), .B(n_1150), .CI(b_mantissa[15]), .CO(n_945), 
      .S(n_944));
   FA_X1 i_473 (.A(n_927), .B(n_925), .CI(n_923), .CO(n_947), .S(n_946));
   FA_X1 i_474 (.A(n_929), .B(n_944), .CI(n_942), .CO(n_949), .S(n_948));
   FA_X1 i_475 (.A(n_940), .B(n_931), .CI(n_946), .CO(n_951), .S(n_950));
   FA_X1 i_476 (.A(n_933), .B(n_948), .CI(n_950), .CO(n_953), .S(n_952));
   FA_X1 i_477 (.A(n_935), .B(n_937), .CI(n_952), .CO(n_955), .S(n_954));
   FA_X1 i_478 (.A(a_mantissa[16]), .B(n_1017), .CI(n_1039), .CO(n_957), 
      .S(n_956));
   FA_X1 i_479 (.A(n_1061), .B(n_1083), .CI(n_1105), .CO(n_959), .S(n_958));
   FA_X1 i_480 (.A(n_1127), .B(b_mantissa[16]), .CI(n_945), .CO(n_961), .S(n_960));
   FA_X1 i_481 (.A(n_943), .B(n_941), .CI(n_947), .CO(n_963), .S(n_962));
   FA_X1 i_482 (.A(n_960), .B(n_958), .CI(n_956), .CO(n_965), .S(n_964));
   FA_X1 i_483 (.A(n_962), .B(n_949), .CI(n_951), .CO(n_967), .S(n_966));
   FA_X1 i_484 (.A(n_964), .B(n_966), .CI(n_953), .CO(n_969), .S(n_968));
   FA_X1 i_485 (.A(a_mantissa[17]), .B(n_1016), .CI(n_1038), .CO(n_971), 
      .S(n_970));
   FA_X1 i_486 (.A(n_1060), .B(n_1082), .CI(n_1104), .CO(n_973), .S(n_972));
   FA_X1 i_487 (.A(b_mantissa[17]), .B(n_959), .CI(n_957), .CO(n_975), .S(n_974));
   FA_X1 i_488 (.A(n_961), .B(n_972), .CI(n_970), .CO(n_977), .S(n_976));
   FA_X1 i_489 (.A(n_963), .B(n_974), .CI(n_965), .CO(n_979), .S(n_978));
   FA_X1 i_490 (.A(n_976), .B(n_967), .CI(n_978), .CO(n_981), .S(n_980));
   FA_X1 i_491 (.A(a_mantissa[18]), .B(n_1015), .CI(n_1037), .CO(n_983), 
      .S(n_982));
   FA_X1 i_492 (.A(n_1059), .B(n_1081), .CI(b_mantissa[18]), .CO(n_985), 
      .S(n_984));
   FA_X1 i_493 (.A(n_973), .B(n_971), .CI(n_975), .CO(n_987), .S(n_986));
   FA_X1 i_494 (.A(n_984), .B(n_982), .CI(n_986), .CO(n_989), .S(n_988));
   FA_X1 i_495 (.A(n_977), .B(n_979), .CI(n_988), .CO(n_991), .S(n_990));
   FA_X1 i_496 (.A(a_mantissa[19]), .B(n_1014), .CI(n_1036), .CO(n_993), 
      .S(n_992));
   FA_X1 i_497 (.A(n_1058), .B(b_mantissa[19]), .CI(n_985), .CO(n_995), .S(n_994));
   FA_X1 i_498 (.A(n_983), .B(n_994), .CI(n_992), .CO(n_997), .S(n_996));
   FA_X1 i_499 (.A(n_987), .B(n_989), .CI(n_996), .CO(n_999), .S(n_998));
   FA_X1 i_500 (.A(a_mantissa[20]), .B(n_1013), .CI(n_1035), .CO(n_1001), 
      .S(n_1000));
   FA_X1 i_501 (.A(b_mantissa[20]), .B(n_993), .CI(n_995), .CO(n_1003), .S(
      n_1002));
   FA_X1 i_502 (.A(n_1000), .B(n_1002), .CI(n_997), .CO(n_1005), .S(n_1004));
   FA_X1 i_503 (.A(a_mantissa[21]), .B(n_1012), .CI(b_mantissa[21]), .CO(n_1007), 
      .S(n_1006));
   FA_X1 i_504 (.A(n_1001), .B(n_1006), .CI(n_1003), .CO(n_1009), .S(n_1008));
   FA_X1 i_505 (.A(a_mantissa[22]), .B(b_mantissa[22]), .CI(n_1007), .CO(n_1011), 
      .S(n_1010));
   NOR2_X1 i_506 (.A1(n_1839), .A2(n_1816), .ZN(n_1012));
   NOR2_X1 i_507 (.A1(n_1839), .A2(n_1815), .ZN(n_1013));
   NOR2_X1 i_508 (.A1(n_1839), .A2(n_1814), .ZN(n_1014));
   NOR2_X1 i_509 (.A1(n_1839), .A2(n_1813), .ZN(n_1015));
   NOR2_X1 i_510 (.A1(n_1839), .A2(n_1812), .ZN(n_1016));
   NOR2_X1 i_511 (.A1(n_1839), .A2(n_1811), .ZN(n_1017));
   NOR2_X1 i_512 (.A1(n_1839), .A2(n_1810), .ZN(n_1018));
   NOR2_X1 i_513 (.A1(n_1839), .A2(n_1809), .ZN(n_1019));
   NOR2_X1 i_514 (.A1(n_1839), .A2(n_1808), .ZN(n_1020));
   NOR2_X1 i_515 (.A1(n_1839), .A2(n_1807), .ZN(n_1021));
   NOR2_X1 i_516 (.A1(n_1839), .A2(n_1806), .ZN(n_1022));
   NOR2_X1 i_517 (.A1(n_1839), .A2(n_1805), .ZN(n_1023));
   NOR2_X1 i_518 (.A1(n_1839), .A2(n_1804), .ZN(n_1024));
   NOR2_X1 i_519 (.A1(n_1839), .A2(n_1803), .ZN(n_1025));
   NOR2_X1 i_520 (.A1(n_1839), .A2(n_1802), .ZN(n_1026));
   NOR2_X1 i_521 (.A1(n_1839), .A2(n_1801), .ZN(n_1027));
   NOR2_X1 i_522 (.A1(n_1839), .A2(n_1800), .ZN(n_1028));
   NOR2_X1 i_523 (.A1(n_1839), .A2(n_1799), .ZN(n_1029));
   NOR2_X1 i_524 (.A1(n_1839), .A2(n_1798), .ZN(n_1030));
   NOR2_X1 i_525 (.A1(n_1839), .A2(n_1797), .ZN(n_1031));
   NOR2_X1 i_526 (.A1(n_1839), .A2(n_1796), .ZN(n_1032));
   NOR2_X1 i_527 (.A1(n_1839), .A2(n_1795), .ZN(n_1033));
   NOR2_X1 i_528 (.A1(n_1839), .A2(n_1794), .ZN(n_1034));
   NOR2_X1 i_529 (.A1(n_1838), .A2(n_1816), .ZN(n_1035));
   NOR2_X1 i_530 (.A1(n_1838), .A2(n_1815), .ZN(n_1036));
   NOR2_X1 i_531 (.A1(n_1838), .A2(n_1814), .ZN(n_1037));
   NOR2_X1 i_532 (.A1(n_1838), .A2(n_1813), .ZN(n_1038));
   NOR2_X1 i_533 (.A1(n_1838), .A2(n_1812), .ZN(n_1039));
   NOR2_X1 i_534 (.A1(n_1838), .A2(n_1811), .ZN(n_1040));
   NOR2_X1 i_535 (.A1(n_1838), .A2(n_1810), .ZN(n_1041));
   NOR2_X1 i_536 (.A1(n_1838), .A2(n_1809), .ZN(n_1042));
   NOR2_X1 i_537 (.A1(n_1838), .A2(n_1808), .ZN(n_1043));
   NOR2_X1 i_538 (.A1(n_1838), .A2(n_1807), .ZN(n_1044));
   NOR2_X1 i_539 (.A1(n_1838), .A2(n_1806), .ZN(n_1045));
   NOR2_X1 i_540 (.A1(n_1838), .A2(n_1805), .ZN(n_1046));
   NOR2_X1 i_541 (.A1(n_1838), .A2(n_1804), .ZN(n_1047));
   NOR2_X1 i_542 (.A1(n_1838), .A2(n_1803), .ZN(n_1048));
   NOR2_X1 i_543 (.A1(n_1838), .A2(n_1802), .ZN(n_1049));
   NOR2_X1 i_544 (.A1(n_1838), .A2(n_1801), .ZN(n_1050));
   NOR2_X1 i_545 (.A1(n_1838), .A2(n_1800), .ZN(n_1051));
   NOR2_X1 i_546 (.A1(n_1838), .A2(n_1799), .ZN(n_1052));
   NOR2_X1 i_547 (.A1(n_1838), .A2(n_1798), .ZN(n_1053));
   NOR2_X1 i_548 (.A1(n_1838), .A2(n_1797), .ZN(n_1054));
   NOR2_X1 i_549 (.A1(n_1838), .A2(n_1796), .ZN(n_1055));
   NOR2_X1 i_550 (.A1(n_1838), .A2(n_1795), .ZN(n_1056));
   NOR2_X1 i_551 (.A1(n_1838), .A2(n_1794), .ZN(n_1057));
   NOR2_X1 i_552 (.A1(n_1837), .A2(n_1816), .ZN(n_1058));
   NOR2_X1 i_553 (.A1(n_1837), .A2(n_1815), .ZN(n_1059));
   NOR2_X1 i_554 (.A1(n_1837), .A2(n_1814), .ZN(n_1060));
   NOR2_X1 i_555 (.A1(n_1837), .A2(n_1813), .ZN(n_1061));
   NOR2_X1 i_556 (.A1(n_1837), .A2(n_1812), .ZN(n_1062));
   NOR2_X1 i_557 (.A1(n_1837), .A2(n_1811), .ZN(n_1063));
   NOR2_X1 i_558 (.A1(n_1837), .A2(n_1810), .ZN(n_1064));
   NOR2_X1 i_559 (.A1(n_1837), .A2(n_1809), .ZN(n_1065));
   NOR2_X1 i_560 (.A1(n_1837), .A2(n_1808), .ZN(n_1066));
   NOR2_X1 i_561 (.A1(n_1837), .A2(n_1807), .ZN(n_1067));
   NOR2_X1 i_562 (.A1(n_1837), .A2(n_1806), .ZN(n_1068));
   NOR2_X1 i_563 (.A1(n_1837), .A2(n_1805), .ZN(n_1069));
   NOR2_X1 i_564 (.A1(n_1837), .A2(n_1804), .ZN(n_1070));
   NOR2_X1 i_565 (.A1(n_1837), .A2(n_1803), .ZN(n_1071));
   NOR2_X1 i_566 (.A1(n_1837), .A2(n_1802), .ZN(n_1072));
   NOR2_X1 i_567 (.A1(n_1837), .A2(n_1801), .ZN(n_1073));
   NOR2_X1 i_568 (.A1(n_1837), .A2(n_1800), .ZN(n_1074));
   NOR2_X1 i_569 (.A1(n_1837), .A2(n_1799), .ZN(n_1075));
   NOR2_X1 i_570 (.A1(n_1837), .A2(n_1798), .ZN(n_1076));
   NOR2_X1 i_571 (.A1(n_1837), .A2(n_1797), .ZN(n_1077));
   NOR2_X1 i_572 (.A1(n_1837), .A2(n_1796), .ZN(n_1078));
   NOR2_X1 i_573 (.A1(n_1837), .A2(n_1795), .ZN(n_1079));
   NOR2_X1 i_574 (.A1(n_1837), .A2(n_1794), .ZN(n_1080));
   NOR2_X1 i_575 (.A1(n_1836), .A2(n_1816), .ZN(n_1081));
   NOR2_X1 i_576 (.A1(n_1836), .A2(n_1815), .ZN(n_1082));
   NOR2_X1 i_577 (.A1(n_1836), .A2(n_1814), .ZN(n_1083));
   NOR2_X1 i_578 (.A1(n_1836), .A2(n_1813), .ZN(n_1084));
   NOR2_X1 i_579 (.A1(n_1836), .A2(n_1812), .ZN(n_1085));
   NOR2_X1 i_580 (.A1(n_1836), .A2(n_1811), .ZN(n_1086));
   NOR2_X1 i_581 (.A1(n_1836), .A2(n_1810), .ZN(n_1087));
   NOR2_X1 i_582 (.A1(n_1836), .A2(n_1809), .ZN(n_1088));
   NOR2_X1 i_583 (.A1(n_1836), .A2(n_1808), .ZN(n_1089));
   NOR2_X1 i_584 (.A1(n_1836), .A2(n_1807), .ZN(n_1090));
   NOR2_X1 i_585 (.A1(n_1836), .A2(n_1806), .ZN(n_1091));
   NOR2_X1 i_586 (.A1(n_1836), .A2(n_1805), .ZN(n_1092));
   NOR2_X1 i_587 (.A1(n_1836), .A2(n_1804), .ZN(n_1093));
   NOR2_X1 i_588 (.A1(n_1836), .A2(n_1803), .ZN(n_1094));
   NOR2_X1 i_589 (.A1(n_1836), .A2(n_1802), .ZN(n_1095));
   NOR2_X1 i_590 (.A1(n_1836), .A2(n_1801), .ZN(n_1096));
   NOR2_X1 i_591 (.A1(n_1836), .A2(n_1800), .ZN(n_1097));
   NOR2_X1 i_592 (.A1(n_1836), .A2(n_1799), .ZN(n_1098));
   NOR2_X1 i_593 (.A1(n_1836), .A2(n_1798), .ZN(n_1099));
   NOR2_X1 i_594 (.A1(n_1836), .A2(n_1797), .ZN(n_1100));
   NOR2_X1 i_595 (.A1(n_1836), .A2(n_1796), .ZN(n_1101));
   NOR2_X1 i_596 (.A1(n_1836), .A2(n_1795), .ZN(n_1102));
   NOR2_X1 i_597 (.A1(n_1836), .A2(n_1794), .ZN(n_1103));
   NOR2_X1 i_598 (.A1(n_1835), .A2(n_1816), .ZN(n_1104));
   NOR2_X1 i_599 (.A1(n_1835), .A2(n_1815), .ZN(n_1105));
   NOR2_X1 i_600 (.A1(n_1835), .A2(n_1814), .ZN(n_1106));
   NOR2_X1 i_601 (.A1(n_1835), .A2(n_1813), .ZN(n_1107));
   NOR2_X1 i_602 (.A1(n_1835), .A2(n_1812), .ZN(n_1108));
   NOR2_X1 i_603 (.A1(n_1835), .A2(n_1811), .ZN(n_1109));
   NOR2_X1 i_604 (.A1(n_1835), .A2(n_1810), .ZN(n_1110));
   NOR2_X1 i_605 (.A1(n_1835), .A2(n_1809), .ZN(n_1111));
   NOR2_X1 i_606 (.A1(n_1835), .A2(n_1808), .ZN(n_1112));
   NOR2_X1 i_607 (.A1(n_1835), .A2(n_1807), .ZN(n_1113));
   NOR2_X1 i_608 (.A1(n_1835), .A2(n_1806), .ZN(n_1114));
   NOR2_X1 i_609 (.A1(n_1835), .A2(n_1805), .ZN(n_1115));
   NOR2_X1 i_610 (.A1(n_1835), .A2(n_1804), .ZN(n_1116));
   NOR2_X1 i_611 (.A1(n_1835), .A2(n_1803), .ZN(n_1117));
   NOR2_X1 i_612 (.A1(n_1835), .A2(n_1802), .ZN(n_1118));
   NOR2_X1 i_613 (.A1(n_1835), .A2(n_1801), .ZN(n_1119));
   NOR2_X1 i_614 (.A1(n_1835), .A2(n_1800), .ZN(n_1120));
   NOR2_X1 i_615 (.A1(n_1835), .A2(n_1799), .ZN(n_1121));
   NOR2_X1 i_616 (.A1(n_1835), .A2(n_1798), .ZN(n_1122));
   NOR2_X1 i_617 (.A1(n_1835), .A2(n_1797), .ZN(n_1123));
   NOR2_X1 i_618 (.A1(n_1835), .A2(n_1796), .ZN(n_1124));
   NOR2_X1 i_619 (.A1(n_1835), .A2(n_1795), .ZN(n_1125));
   NOR2_X1 i_620 (.A1(n_1835), .A2(n_1794), .ZN(n_1126));
   NOR2_X1 i_621 (.A1(n_1834), .A2(n_1816), .ZN(n_1127));
   NOR2_X1 i_622 (.A1(n_1834), .A2(n_1815), .ZN(n_1128));
   NOR2_X1 i_623 (.A1(n_1834), .A2(n_1814), .ZN(n_1129));
   NOR2_X1 i_624 (.A1(n_1834), .A2(n_1813), .ZN(n_1130));
   NOR2_X1 i_625 (.A1(n_1834), .A2(n_1812), .ZN(n_1131));
   NOR2_X1 i_626 (.A1(n_1834), .A2(n_1811), .ZN(n_1132));
   NOR2_X1 i_627 (.A1(n_1834), .A2(n_1810), .ZN(n_1133));
   NOR2_X1 i_628 (.A1(n_1834), .A2(n_1809), .ZN(n_1134));
   NOR2_X1 i_629 (.A1(n_1834), .A2(n_1808), .ZN(n_1135));
   NOR2_X1 i_630 (.A1(n_1834), .A2(n_1807), .ZN(n_1136));
   NOR2_X1 i_631 (.A1(n_1834), .A2(n_1806), .ZN(n_1137));
   NOR2_X1 i_632 (.A1(n_1834), .A2(n_1805), .ZN(n_1138));
   NOR2_X1 i_633 (.A1(n_1834), .A2(n_1804), .ZN(n_1139));
   NOR2_X1 i_634 (.A1(n_1834), .A2(n_1803), .ZN(n_1140));
   NOR2_X1 i_635 (.A1(n_1834), .A2(n_1802), .ZN(n_1141));
   NOR2_X1 i_636 (.A1(n_1834), .A2(n_1801), .ZN(n_1142));
   NOR2_X1 i_637 (.A1(n_1834), .A2(n_1800), .ZN(n_1143));
   NOR2_X1 i_638 (.A1(n_1834), .A2(n_1799), .ZN(n_1144));
   NOR2_X1 i_639 (.A1(n_1834), .A2(n_1798), .ZN(n_1145));
   NOR2_X1 i_640 (.A1(n_1834), .A2(n_1797), .ZN(n_1146));
   NOR2_X1 i_641 (.A1(n_1834), .A2(n_1796), .ZN(n_1147));
   NOR2_X1 i_642 (.A1(n_1834), .A2(n_1795), .ZN(n_1148));
   NOR2_X1 i_643 (.A1(n_1834), .A2(n_1794), .ZN(n_1149));
   NOR2_X1 i_644 (.A1(n_1833), .A2(n_1816), .ZN(n_1150));
   NOR2_X1 i_645 (.A1(n_1833), .A2(n_1815), .ZN(n_1151));
   NOR2_X1 i_646 (.A1(n_1833), .A2(n_1814), .ZN(n_1152));
   NOR2_X1 i_647 (.A1(n_1833), .A2(n_1813), .ZN(n_1153));
   NOR2_X1 i_648 (.A1(n_1833), .A2(n_1812), .ZN(n_1154));
   NOR2_X1 i_649 (.A1(n_1833), .A2(n_1811), .ZN(n_1155));
   NOR2_X1 i_650 (.A1(n_1833), .A2(n_1810), .ZN(n_1156));
   NOR2_X1 i_651 (.A1(n_1833), .A2(n_1809), .ZN(n_1157));
   NOR2_X1 i_652 (.A1(n_1833), .A2(n_1808), .ZN(n_1158));
   NOR2_X1 i_653 (.A1(n_1833), .A2(n_1807), .ZN(n_1159));
   NOR2_X1 i_654 (.A1(n_1833), .A2(n_1806), .ZN(n_1160));
   NOR2_X1 i_655 (.A1(n_1833), .A2(n_1805), .ZN(n_1161));
   NOR2_X1 i_656 (.A1(n_1833), .A2(n_1804), .ZN(n_1162));
   NOR2_X1 i_657 (.A1(n_1833), .A2(n_1803), .ZN(n_1163));
   NOR2_X1 i_658 (.A1(n_1833), .A2(n_1802), .ZN(n_1164));
   NOR2_X1 i_659 (.A1(n_1833), .A2(n_1801), .ZN(n_1165));
   NOR2_X1 i_660 (.A1(n_1833), .A2(n_1800), .ZN(n_1166));
   NOR2_X1 i_661 (.A1(n_1833), .A2(n_1799), .ZN(n_1167));
   NOR2_X1 i_662 (.A1(n_1833), .A2(n_1798), .ZN(n_1168));
   NOR2_X1 i_663 (.A1(n_1833), .A2(n_1797), .ZN(n_1169));
   NOR2_X1 i_664 (.A1(n_1833), .A2(n_1796), .ZN(n_1170));
   NOR2_X1 i_665 (.A1(n_1833), .A2(n_1795), .ZN(n_1171));
   NOR2_X1 i_666 (.A1(n_1833), .A2(n_1794), .ZN(n_1172));
   NOR2_X1 i_667 (.A1(n_1832), .A2(n_1816), .ZN(n_1173));
   NOR2_X1 i_668 (.A1(n_1832), .A2(n_1815), .ZN(n_1174));
   NOR2_X1 i_669 (.A1(n_1832), .A2(n_1814), .ZN(n_1175));
   NOR2_X1 i_670 (.A1(n_1832), .A2(n_1813), .ZN(n_1176));
   NOR2_X1 i_671 (.A1(n_1832), .A2(n_1812), .ZN(n_1177));
   NOR2_X1 i_672 (.A1(n_1832), .A2(n_1811), .ZN(n_1178));
   NOR2_X1 i_673 (.A1(n_1832), .A2(n_1810), .ZN(n_1179));
   NOR2_X1 i_674 (.A1(n_1832), .A2(n_1809), .ZN(n_1180));
   NOR2_X1 i_675 (.A1(n_1832), .A2(n_1808), .ZN(n_1181));
   NOR2_X1 i_676 (.A1(n_1832), .A2(n_1807), .ZN(n_1182));
   NOR2_X1 i_677 (.A1(n_1832), .A2(n_1806), .ZN(n_1183));
   NOR2_X1 i_678 (.A1(n_1832), .A2(n_1805), .ZN(n_1184));
   NOR2_X1 i_679 (.A1(n_1832), .A2(n_1804), .ZN(n_1185));
   NOR2_X1 i_680 (.A1(n_1832), .A2(n_1803), .ZN(n_1186));
   NOR2_X1 i_681 (.A1(n_1832), .A2(n_1802), .ZN(n_1187));
   NOR2_X1 i_682 (.A1(n_1832), .A2(n_1801), .ZN(n_1188));
   NOR2_X1 i_683 (.A1(n_1832), .A2(n_1800), .ZN(n_1189));
   NOR2_X1 i_684 (.A1(n_1832), .A2(n_1799), .ZN(n_1190));
   NOR2_X1 i_685 (.A1(n_1832), .A2(n_1798), .ZN(n_1191));
   NOR2_X1 i_686 (.A1(n_1832), .A2(n_1797), .ZN(n_1192));
   NOR2_X1 i_687 (.A1(n_1832), .A2(n_1796), .ZN(n_1193));
   NOR2_X1 i_688 (.A1(n_1832), .A2(n_1795), .ZN(n_1194));
   NOR2_X1 i_689 (.A1(n_1832), .A2(n_1794), .ZN(n_1195));
   NOR2_X1 i_690 (.A1(n_1831), .A2(n_1816), .ZN(n_1196));
   NOR2_X1 i_691 (.A1(n_1831), .A2(n_1815), .ZN(n_1197));
   NOR2_X1 i_692 (.A1(n_1831), .A2(n_1814), .ZN(n_1198));
   NOR2_X1 i_693 (.A1(n_1831), .A2(n_1813), .ZN(n_1199));
   NOR2_X1 i_694 (.A1(n_1831), .A2(n_1812), .ZN(n_1200));
   NOR2_X1 i_695 (.A1(n_1831), .A2(n_1811), .ZN(n_1201));
   NOR2_X1 i_696 (.A1(n_1831), .A2(n_1810), .ZN(n_1202));
   NOR2_X1 i_697 (.A1(n_1831), .A2(n_1809), .ZN(n_1203));
   NOR2_X1 i_698 (.A1(n_1831), .A2(n_1808), .ZN(n_1204));
   NOR2_X1 i_699 (.A1(n_1831), .A2(n_1807), .ZN(n_1205));
   NOR2_X1 i_700 (.A1(n_1831), .A2(n_1806), .ZN(n_1206));
   NOR2_X1 i_701 (.A1(n_1831), .A2(n_1805), .ZN(n_1207));
   NOR2_X1 i_702 (.A1(n_1831), .A2(n_1804), .ZN(n_1208));
   NOR2_X1 i_703 (.A1(n_1831), .A2(n_1803), .ZN(n_1209));
   NOR2_X1 i_704 (.A1(n_1831), .A2(n_1802), .ZN(n_1210));
   NOR2_X1 i_705 (.A1(n_1831), .A2(n_1801), .ZN(n_1211));
   NOR2_X1 i_706 (.A1(n_1831), .A2(n_1800), .ZN(n_1212));
   NOR2_X1 i_707 (.A1(n_1831), .A2(n_1799), .ZN(n_1213));
   NOR2_X1 i_708 (.A1(n_1831), .A2(n_1798), .ZN(n_1214));
   NOR2_X1 i_709 (.A1(n_1831), .A2(n_1797), .ZN(n_1215));
   NOR2_X1 i_710 (.A1(n_1831), .A2(n_1796), .ZN(n_1216));
   NOR2_X1 i_711 (.A1(n_1831), .A2(n_1795), .ZN(n_1217));
   NOR2_X1 i_712 (.A1(n_1831), .A2(n_1794), .ZN(n_1218));
   NOR2_X1 i_713 (.A1(n_1830), .A2(n_1816), .ZN(n_1219));
   NOR2_X1 i_714 (.A1(n_1830), .A2(n_1815), .ZN(n_1220));
   NOR2_X1 i_715 (.A1(n_1830), .A2(n_1814), .ZN(n_1221));
   NOR2_X1 i_716 (.A1(n_1830), .A2(n_1813), .ZN(n_1222));
   NOR2_X1 i_717 (.A1(n_1830), .A2(n_1812), .ZN(n_1223));
   NOR2_X1 i_718 (.A1(n_1830), .A2(n_1811), .ZN(n_1224));
   NOR2_X1 i_719 (.A1(n_1830), .A2(n_1810), .ZN(n_1225));
   NOR2_X1 i_720 (.A1(n_1830), .A2(n_1809), .ZN(n_1226));
   NOR2_X1 i_721 (.A1(n_1830), .A2(n_1808), .ZN(n_1227));
   NOR2_X1 i_722 (.A1(n_1830), .A2(n_1807), .ZN(n_1228));
   NOR2_X1 i_723 (.A1(n_1830), .A2(n_1806), .ZN(n_1229));
   NOR2_X1 i_724 (.A1(n_1830), .A2(n_1805), .ZN(n_1230));
   NOR2_X1 i_725 (.A1(n_1830), .A2(n_1804), .ZN(n_1231));
   NOR2_X1 i_726 (.A1(n_1830), .A2(n_1803), .ZN(n_1232));
   NOR2_X1 i_727 (.A1(n_1830), .A2(n_1802), .ZN(n_1233));
   NOR2_X1 i_728 (.A1(n_1830), .A2(n_1801), .ZN(n_1234));
   NOR2_X1 i_729 (.A1(n_1830), .A2(n_1800), .ZN(n_1235));
   NOR2_X1 i_730 (.A1(n_1830), .A2(n_1799), .ZN(n_1236));
   NOR2_X1 i_731 (.A1(n_1830), .A2(n_1798), .ZN(n_1237));
   NOR2_X1 i_732 (.A1(n_1830), .A2(n_1797), .ZN(n_1238));
   NOR2_X1 i_733 (.A1(n_1830), .A2(n_1796), .ZN(n_1239));
   NOR2_X1 i_734 (.A1(n_1830), .A2(n_1795), .ZN(n_1240));
   NOR2_X1 i_735 (.A1(n_1830), .A2(n_1794), .ZN(n_1241));
   NOR2_X1 i_736 (.A1(n_1829), .A2(n_1816), .ZN(n_1242));
   NOR2_X1 i_737 (.A1(n_1829), .A2(n_1815), .ZN(n_1243));
   NOR2_X1 i_738 (.A1(n_1829), .A2(n_1814), .ZN(n_1244));
   NOR2_X1 i_739 (.A1(n_1829), .A2(n_1813), .ZN(n_1245));
   NOR2_X1 i_740 (.A1(n_1829), .A2(n_1812), .ZN(n_1246));
   NOR2_X1 i_741 (.A1(n_1829), .A2(n_1811), .ZN(n_1247));
   NOR2_X1 i_742 (.A1(n_1829), .A2(n_1810), .ZN(n_1248));
   NOR2_X1 i_743 (.A1(n_1829), .A2(n_1809), .ZN(n_1249));
   NOR2_X1 i_744 (.A1(n_1829), .A2(n_1808), .ZN(n_1250));
   NOR2_X1 i_745 (.A1(n_1829), .A2(n_1807), .ZN(n_1251));
   NOR2_X1 i_746 (.A1(n_1829), .A2(n_1806), .ZN(n_1252));
   NOR2_X1 i_747 (.A1(n_1829), .A2(n_1805), .ZN(n_1253));
   NOR2_X1 i_748 (.A1(n_1829), .A2(n_1804), .ZN(n_1254));
   NOR2_X1 i_749 (.A1(n_1829), .A2(n_1803), .ZN(n_1255));
   NOR2_X1 i_750 (.A1(n_1829), .A2(n_1802), .ZN(n_1256));
   NOR2_X1 i_751 (.A1(n_1829), .A2(n_1801), .ZN(n_1257));
   NOR2_X1 i_752 (.A1(n_1829), .A2(n_1800), .ZN(n_1258));
   NOR2_X1 i_753 (.A1(n_1829), .A2(n_1799), .ZN(n_1259));
   NOR2_X1 i_754 (.A1(n_1829), .A2(n_1798), .ZN(n_1260));
   NOR2_X1 i_755 (.A1(n_1829), .A2(n_1797), .ZN(n_1261));
   NOR2_X1 i_756 (.A1(n_1829), .A2(n_1796), .ZN(n_1262));
   NOR2_X1 i_757 (.A1(n_1829), .A2(n_1795), .ZN(n_1263));
   NOR2_X1 i_758 (.A1(n_1829), .A2(n_1794), .ZN(n_1264));
   NOR2_X1 i_759 (.A1(n_1828), .A2(n_1816), .ZN(n_1265));
   NOR2_X1 i_760 (.A1(n_1828), .A2(n_1815), .ZN(n_1266));
   NOR2_X1 i_761 (.A1(n_1828), .A2(n_1814), .ZN(n_1267));
   NOR2_X1 i_762 (.A1(n_1828), .A2(n_1813), .ZN(n_1268));
   NOR2_X1 i_763 (.A1(n_1828), .A2(n_1812), .ZN(n_1269));
   NOR2_X1 i_764 (.A1(n_1828), .A2(n_1811), .ZN(n_1270));
   NOR2_X1 i_765 (.A1(n_1828), .A2(n_1810), .ZN(n_1271));
   NOR2_X1 i_766 (.A1(n_1828), .A2(n_1809), .ZN(n_1272));
   NOR2_X1 i_767 (.A1(n_1828), .A2(n_1808), .ZN(n_1273));
   NOR2_X1 i_768 (.A1(n_1828), .A2(n_1807), .ZN(n_1274));
   NOR2_X1 i_769 (.A1(n_1828), .A2(n_1806), .ZN(n_1275));
   NOR2_X1 i_770 (.A1(n_1828), .A2(n_1805), .ZN(n_1276));
   NOR2_X1 i_771 (.A1(n_1828), .A2(n_1804), .ZN(n_1277));
   NOR2_X1 i_772 (.A1(n_1828), .A2(n_1803), .ZN(n_1278));
   NOR2_X1 i_773 (.A1(n_1828), .A2(n_1802), .ZN(n_1279));
   NOR2_X1 i_774 (.A1(n_1828), .A2(n_1801), .ZN(n_1280));
   NOR2_X1 i_775 (.A1(n_1828), .A2(n_1800), .ZN(n_1281));
   NOR2_X1 i_776 (.A1(n_1828), .A2(n_1799), .ZN(n_1282));
   NOR2_X1 i_777 (.A1(n_1828), .A2(n_1798), .ZN(n_1283));
   NOR2_X1 i_778 (.A1(n_1828), .A2(n_1797), .ZN(n_1284));
   NOR2_X1 i_779 (.A1(n_1828), .A2(n_1796), .ZN(n_1285));
   NOR2_X1 i_780 (.A1(n_1828), .A2(n_1795), .ZN(n_1286));
   NOR2_X1 i_781 (.A1(n_1828), .A2(n_1794), .ZN(n_1287));
   NOR2_X1 i_782 (.A1(n_1827), .A2(n_1816), .ZN(n_1288));
   NOR2_X1 i_783 (.A1(n_1827), .A2(n_1815), .ZN(n_1289));
   NOR2_X1 i_784 (.A1(n_1827), .A2(n_1814), .ZN(n_1290));
   NOR2_X1 i_785 (.A1(n_1827), .A2(n_1813), .ZN(n_1291));
   NOR2_X1 i_786 (.A1(n_1827), .A2(n_1812), .ZN(n_1292));
   NOR2_X1 i_787 (.A1(n_1827), .A2(n_1811), .ZN(n_1293));
   NOR2_X1 i_788 (.A1(n_1827), .A2(n_1810), .ZN(n_1294));
   NOR2_X1 i_789 (.A1(n_1827), .A2(n_1809), .ZN(n_1295));
   NOR2_X1 i_790 (.A1(n_1827), .A2(n_1808), .ZN(n_1296));
   NOR2_X1 i_791 (.A1(n_1827), .A2(n_1807), .ZN(n_1297));
   NOR2_X1 i_792 (.A1(n_1827), .A2(n_1806), .ZN(n_1298));
   NOR2_X1 i_793 (.A1(n_1827), .A2(n_1805), .ZN(n_1299));
   NOR2_X1 i_794 (.A1(n_1827), .A2(n_1804), .ZN(n_1300));
   NOR2_X1 i_795 (.A1(n_1827), .A2(n_1803), .ZN(n_1301));
   NOR2_X1 i_796 (.A1(n_1827), .A2(n_1802), .ZN(n_1302));
   NOR2_X1 i_797 (.A1(n_1827), .A2(n_1801), .ZN(n_1303));
   NOR2_X1 i_798 (.A1(n_1827), .A2(n_1800), .ZN(n_1304));
   NOR2_X1 i_799 (.A1(n_1827), .A2(n_1799), .ZN(n_1305));
   NOR2_X1 i_800 (.A1(n_1827), .A2(n_1798), .ZN(n_1306));
   NOR2_X1 i_801 (.A1(n_1827), .A2(n_1797), .ZN(n_1307));
   NOR2_X1 i_802 (.A1(n_1827), .A2(n_1796), .ZN(n_1308));
   NOR2_X1 i_803 (.A1(n_1827), .A2(n_1795), .ZN(n_1309));
   NOR2_X1 i_804 (.A1(n_1827), .A2(n_1794), .ZN(n_1310));
   NOR2_X1 i_805 (.A1(n_1826), .A2(n_1816), .ZN(n_1311));
   NOR2_X1 i_806 (.A1(n_1826), .A2(n_1815), .ZN(n_1312));
   NOR2_X1 i_807 (.A1(n_1826), .A2(n_1814), .ZN(n_1313));
   NOR2_X1 i_808 (.A1(n_1826), .A2(n_1813), .ZN(n_1314));
   NOR2_X1 i_809 (.A1(n_1826), .A2(n_1812), .ZN(n_1315));
   NOR2_X1 i_810 (.A1(n_1826), .A2(n_1811), .ZN(n_1316));
   NOR2_X1 i_811 (.A1(n_1826), .A2(n_1810), .ZN(n_1317));
   NOR2_X1 i_812 (.A1(n_1826), .A2(n_1809), .ZN(n_1318));
   NOR2_X1 i_813 (.A1(n_1826), .A2(n_1808), .ZN(n_1319));
   NOR2_X1 i_814 (.A1(n_1826), .A2(n_1807), .ZN(n_1320));
   NOR2_X1 i_815 (.A1(n_1826), .A2(n_1806), .ZN(n_1321));
   NOR2_X1 i_816 (.A1(n_1826), .A2(n_1805), .ZN(n_1322));
   NOR2_X1 i_817 (.A1(n_1826), .A2(n_1804), .ZN(n_1323));
   NOR2_X1 i_818 (.A1(n_1826), .A2(n_1803), .ZN(n_1324));
   NOR2_X1 i_819 (.A1(n_1826), .A2(n_1802), .ZN(n_1325));
   NOR2_X1 i_820 (.A1(n_1826), .A2(n_1801), .ZN(n_1326));
   NOR2_X1 i_821 (.A1(n_1826), .A2(n_1800), .ZN(n_1327));
   NOR2_X1 i_822 (.A1(n_1826), .A2(n_1799), .ZN(n_1328));
   NOR2_X1 i_823 (.A1(n_1826), .A2(n_1798), .ZN(n_1329));
   NOR2_X1 i_824 (.A1(n_1826), .A2(n_1797), .ZN(n_1330));
   NOR2_X1 i_825 (.A1(n_1826), .A2(n_1796), .ZN(n_1331));
   NOR2_X1 i_826 (.A1(n_1826), .A2(n_1795), .ZN(n_1332));
   NOR2_X1 i_827 (.A1(n_1826), .A2(n_1794), .ZN(n_1333));
   NOR2_X1 i_828 (.A1(n_1825), .A2(n_1816), .ZN(n_1334));
   NOR2_X1 i_829 (.A1(n_1825), .A2(n_1815), .ZN(n_1335));
   NOR2_X1 i_830 (.A1(n_1825), .A2(n_1814), .ZN(n_1336));
   NOR2_X1 i_831 (.A1(n_1825), .A2(n_1813), .ZN(n_1337));
   NOR2_X1 i_832 (.A1(n_1825), .A2(n_1812), .ZN(n_1338));
   NOR2_X1 i_833 (.A1(n_1825), .A2(n_1811), .ZN(n_1339));
   NOR2_X1 i_834 (.A1(n_1825), .A2(n_1810), .ZN(n_1340));
   NOR2_X1 i_835 (.A1(n_1825), .A2(n_1809), .ZN(n_1341));
   NOR2_X1 i_836 (.A1(n_1825), .A2(n_1808), .ZN(n_1342));
   NOR2_X1 i_837 (.A1(n_1825), .A2(n_1807), .ZN(n_1343));
   NOR2_X1 i_838 (.A1(n_1825), .A2(n_1806), .ZN(n_1344));
   NOR2_X1 i_839 (.A1(n_1825), .A2(n_1805), .ZN(n_1345));
   NOR2_X1 i_840 (.A1(n_1825), .A2(n_1804), .ZN(n_1346));
   NOR2_X1 i_841 (.A1(n_1825), .A2(n_1803), .ZN(n_1347));
   NOR2_X1 i_842 (.A1(n_1825), .A2(n_1802), .ZN(n_1348));
   NOR2_X1 i_843 (.A1(n_1825), .A2(n_1801), .ZN(n_1349));
   NOR2_X1 i_844 (.A1(n_1825), .A2(n_1800), .ZN(n_1350));
   NOR2_X1 i_845 (.A1(n_1825), .A2(n_1799), .ZN(n_1351));
   NOR2_X1 i_846 (.A1(n_1825), .A2(n_1798), .ZN(n_1352));
   NOR2_X1 i_847 (.A1(n_1825), .A2(n_1797), .ZN(n_1353));
   NOR2_X1 i_848 (.A1(n_1825), .A2(n_1796), .ZN(n_1354));
   NOR2_X1 i_849 (.A1(n_1825), .A2(n_1795), .ZN(n_1355));
   NOR2_X1 i_850 (.A1(n_1825), .A2(n_1794), .ZN(n_1356));
   NOR2_X1 i_851 (.A1(n_1824), .A2(n_1816), .ZN(n_1357));
   NOR2_X1 i_852 (.A1(n_1824), .A2(n_1815), .ZN(n_1358));
   NOR2_X1 i_853 (.A1(n_1824), .A2(n_1814), .ZN(n_1359));
   NOR2_X1 i_854 (.A1(n_1824), .A2(n_1813), .ZN(n_1360));
   NOR2_X1 i_855 (.A1(n_1824), .A2(n_1812), .ZN(n_1361));
   NOR2_X1 i_856 (.A1(n_1824), .A2(n_1811), .ZN(n_1362));
   NOR2_X1 i_857 (.A1(n_1824), .A2(n_1810), .ZN(n_1363));
   NOR2_X1 i_858 (.A1(n_1824), .A2(n_1809), .ZN(n_1364));
   NOR2_X1 i_859 (.A1(n_1824), .A2(n_1808), .ZN(n_1365));
   NOR2_X1 i_860 (.A1(n_1824), .A2(n_1807), .ZN(n_1366));
   NOR2_X1 i_861 (.A1(n_1824), .A2(n_1806), .ZN(n_1367));
   NOR2_X1 i_862 (.A1(n_1824), .A2(n_1805), .ZN(n_1368));
   NOR2_X1 i_863 (.A1(n_1824), .A2(n_1804), .ZN(n_1369));
   NOR2_X1 i_864 (.A1(n_1824), .A2(n_1803), .ZN(n_1370));
   NOR2_X1 i_865 (.A1(n_1824), .A2(n_1802), .ZN(n_1371));
   NOR2_X1 i_866 (.A1(n_1824), .A2(n_1801), .ZN(n_1372));
   NOR2_X1 i_867 (.A1(n_1824), .A2(n_1800), .ZN(n_1373));
   NOR2_X1 i_868 (.A1(n_1824), .A2(n_1799), .ZN(n_1374));
   NOR2_X1 i_869 (.A1(n_1824), .A2(n_1798), .ZN(n_1375));
   NOR2_X1 i_870 (.A1(n_1824), .A2(n_1797), .ZN(n_1376));
   NOR2_X1 i_871 (.A1(n_1824), .A2(n_1796), .ZN(n_1377));
   NOR2_X1 i_872 (.A1(n_1824), .A2(n_1795), .ZN(n_1378));
   NOR2_X1 i_873 (.A1(n_1824), .A2(n_1794), .ZN(n_1379));
   NOR2_X1 i_874 (.A1(n_1823), .A2(n_1816), .ZN(n_1380));
   NOR2_X1 i_875 (.A1(n_1823), .A2(n_1815), .ZN(n_1381));
   NOR2_X1 i_876 (.A1(n_1823), .A2(n_1814), .ZN(n_1382));
   NOR2_X1 i_877 (.A1(n_1823), .A2(n_1813), .ZN(n_1383));
   NOR2_X1 i_878 (.A1(n_1823), .A2(n_1812), .ZN(n_1384));
   NOR2_X1 i_879 (.A1(n_1823), .A2(n_1811), .ZN(n_1385));
   NOR2_X1 i_880 (.A1(n_1823), .A2(n_1810), .ZN(n_1386));
   NOR2_X1 i_881 (.A1(n_1823), .A2(n_1809), .ZN(n_1387));
   NOR2_X1 i_882 (.A1(n_1823), .A2(n_1808), .ZN(n_1388));
   NOR2_X1 i_883 (.A1(n_1823), .A2(n_1807), .ZN(n_1389));
   NOR2_X1 i_884 (.A1(n_1823), .A2(n_1806), .ZN(n_1390));
   NOR2_X1 i_885 (.A1(n_1823), .A2(n_1805), .ZN(n_1391));
   NOR2_X1 i_886 (.A1(n_1823), .A2(n_1804), .ZN(n_1392));
   NOR2_X1 i_887 (.A1(n_1823), .A2(n_1803), .ZN(n_1393));
   NOR2_X1 i_888 (.A1(n_1823), .A2(n_1802), .ZN(n_1394));
   NOR2_X1 i_889 (.A1(n_1823), .A2(n_1801), .ZN(n_1395));
   NOR2_X1 i_890 (.A1(n_1823), .A2(n_1800), .ZN(n_1396));
   NOR2_X1 i_891 (.A1(n_1823), .A2(n_1799), .ZN(n_1397));
   NOR2_X1 i_892 (.A1(n_1823), .A2(n_1798), .ZN(n_1398));
   NOR2_X1 i_893 (.A1(n_1823), .A2(n_1797), .ZN(n_1399));
   NOR2_X1 i_894 (.A1(n_1823), .A2(n_1796), .ZN(n_1400));
   NOR2_X1 i_895 (.A1(n_1823), .A2(n_1795), .ZN(n_1401));
   NOR2_X1 i_896 (.A1(n_1823), .A2(n_1794), .ZN(n_1402));
   NOR2_X1 i_897 (.A1(n_1822), .A2(n_1816), .ZN(n_1403));
   NOR2_X1 i_898 (.A1(n_1822), .A2(n_1815), .ZN(n_1404));
   NOR2_X1 i_899 (.A1(n_1822), .A2(n_1814), .ZN(n_1405));
   NOR2_X1 i_900 (.A1(n_1822), .A2(n_1813), .ZN(n_1406));
   NOR2_X1 i_901 (.A1(n_1822), .A2(n_1812), .ZN(n_1407));
   NOR2_X1 i_902 (.A1(n_1822), .A2(n_1811), .ZN(n_1408));
   NOR2_X1 i_903 (.A1(n_1822), .A2(n_1810), .ZN(n_1409));
   NOR2_X1 i_904 (.A1(n_1822), .A2(n_1809), .ZN(n_1410));
   NOR2_X1 i_905 (.A1(n_1822), .A2(n_1808), .ZN(n_1411));
   NOR2_X1 i_906 (.A1(n_1822), .A2(n_1807), .ZN(n_1412));
   NOR2_X1 i_907 (.A1(n_1822), .A2(n_1806), .ZN(n_1413));
   NOR2_X1 i_908 (.A1(n_1822), .A2(n_1805), .ZN(n_1414));
   NOR2_X1 i_909 (.A1(n_1822), .A2(n_1804), .ZN(n_1415));
   NOR2_X1 i_910 (.A1(n_1822), .A2(n_1803), .ZN(n_1416));
   NOR2_X1 i_911 (.A1(n_1822), .A2(n_1802), .ZN(n_1417));
   NOR2_X1 i_912 (.A1(n_1822), .A2(n_1801), .ZN(n_1418));
   NOR2_X1 i_913 (.A1(n_1822), .A2(n_1800), .ZN(n_1419));
   NOR2_X1 i_914 (.A1(n_1822), .A2(n_1799), .ZN(n_1420));
   NOR2_X1 i_915 (.A1(n_1822), .A2(n_1798), .ZN(n_1421));
   NOR2_X1 i_916 (.A1(n_1822), .A2(n_1797), .ZN(n_1422));
   NOR2_X1 i_917 (.A1(n_1822), .A2(n_1796), .ZN(n_1423));
   NOR2_X1 i_918 (.A1(n_1822), .A2(n_1795), .ZN(n_1424));
   NOR2_X1 i_919 (.A1(n_1822), .A2(n_1794), .ZN(n_1425));
   NOR2_X1 i_920 (.A1(n_1821), .A2(n_1816), .ZN(n_1426));
   NOR2_X1 i_921 (.A1(n_1821), .A2(n_1815), .ZN(n_1427));
   NOR2_X1 i_922 (.A1(n_1821), .A2(n_1814), .ZN(n_1428));
   NOR2_X1 i_923 (.A1(n_1821), .A2(n_1813), .ZN(n_1429));
   NOR2_X1 i_924 (.A1(n_1821), .A2(n_1812), .ZN(n_1430));
   NOR2_X1 i_925 (.A1(n_1821), .A2(n_1811), .ZN(n_1431));
   NOR2_X1 i_926 (.A1(n_1821), .A2(n_1810), .ZN(n_1432));
   NOR2_X1 i_927 (.A1(n_1821), .A2(n_1809), .ZN(n_1433));
   NOR2_X1 i_928 (.A1(n_1821), .A2(n_1808), .ZN(n_1434));
   NOR2_X1 i_929 (.A1(n_1821), .A2(n_1807), .ZN(n_1435));
   NOR2_X1 i_930 (.A1(n_1821), .A2(n_1806), .ZN(n_1436));
   NOR2_X1 i_931 (.A1(n_1821), .A2(n_1805), .ZN(n_1437));
   NOR2_X1 i_932 (.A1(n_1821), .A2(n_1804), .ZN(n_1438));
   NOR2_X1 i_933 (.A1(n_1821), .A2(n_1803), .ZN(n_1439));
   NOR2_X1 i_934 (.A1(n_1821), .A2(n_1802), .ZN(n_1440));
   NOR2_X1 i_935 (.A1(n_1821), .A2(n_1801), .ZN(n_1441));
   NOR2_X1 i_936 (.A1(n_1821), .A2(n_1800), .ZN(n_1442));
   NOR2_X1 i_937 (.A1(n_1821), .A2(n_1799), .ZN(n_1443));
   NOR2_X1 i_938 (.A1(n_1821), .A2(n_1798), .ZN(n_1444));
   NOR2_X1 i_939 (.A1(n_1821), .A2(n_1797), .ZN(n_1445));
   NOR2_X1 i_940 (.A1(n_1821), .A2(n_1796), .ZN(n_1446));
   NOR2_X1 i_941 (.A1(n_1821), .A2(n_1795), .ZN(n_1447));
   NOR2_X1 i_942 (.A1(n_1821), .A2(n_1794), .ZN(n_1448));
   NOR2_X1 i_943 (.A1(n_1820), .A2(n_1816), .ZN(n_1449));
   NOR2_X1 i_944 (.A1(n_1820), .A2(n_1815), .ZN(n_1450));
   NOR2_X1 i_945 (.A1(n_1820), .A2(n_1814), .ZN(n_1451));
   NOR2_X1 i_946 (.A1(n_1820), .A2(n_1813), .ZN(n_1452));
   NOR2_X1 i_947 (.A1(n_1820), .A2(n_1812), .ZN(n_1453));
   NOR2_X1 i_948 (.A1(n_1820), .A2(n_1811), .ZN(n_1454));
   NOR2_X1 i_949 (.A1(n_1820), .A2(n_1810), .ZN(n_1455));
   NOR2_X1 i_950 (.A1(n_1820), .A2(n_1809), .ZN(n_1456));
   NOR2_X1 i_951 (.A1(n_1820), .A2(n_1808), .ZN(n_1457));
   NOR2_X1 i_952 (.A1(n_1820), .A2(n_1807), .ZN(n_1458));
   NOR2_X1 i_953 (.A1(n_1820), .A2(n_1806), .ZN(n_1459));
   NOR2_X1 i_954 (.A1(n_1820), .A2(n_1805), .ZN(n_1460));
   NOR2_X1 i_955 (.A1(n_1820), .A2(n_1804), .ZN(n_1461));
   NOR2_X1 i_956 (.A1(n_1820), .A2(n_1803), .ZN(n_1462));
   NOR2_X1 i_957 (.A1(n_1820), .A2(n_1802), .ZN(n_1463));
   NOR2_X1 i_958 (.A1(n_1820), .A2(n_1801), .ZN(n_1464));
   NOR2_X1 i_959 (.A1(n_1820), .A2(n_1800), .ZN(n_1465));
   NOR2_X1 i_960 (.A1(n_1820), .A2(n_1799), .ZN(n_1466));
   NOR2_X1 i_961 (.A1(n_1820), .A2(n_1798), .ZN(n_1467));
   NOR2_X1 i_962 (.A1(n_1820), .A2(n_1797), .ZN(n_1468));
   NOR2_X1 i_963 (.A1(n_1820), .A2(n_1796), .ZN(n_1469));
   NOR2_X1 i_964 (.A1(n_1820), .A2(n_1795), .ZN(n_1470));
   NOR2_X1 i_965 (.A1(n_1820), .A2(n_1794), .ZN(n_1471));
   NOR2_X1 i_966 (.A1(n_1819), .A2(n_1816), .ZN(n_1472));
   NOR2_X1 i_967 (.A1(n_1819), .A2(n_1815), .ZN(n_1473));
   NOR2_X1 i_968 (.A1(n_1819), .A2(n_1814), .ZN(n_1474));
   NOR2_X1 i_969 (.A1(n_1819), .A2(n_1813), .ZN(n_1475));
   NOR2_X1 i_970 (.A1(n_1819), .A2(n_1812), .ZN(n_1476));
   NOR2_X1 i_971 (.A1(n_1819), .A2(n_1811), .ZN(n_1477));
   NOR2_X1 i_972 (.A1(n_1819), .A2(n_1810), .ZN(n_1478));
   NOR2_X1 i_973 (.A1(n_1819), .A2(n_1809), .ZN(n_1479));
   NOR2_X1 i_974 (.A1(n_1819), .A2(n_1808), .ZN(n_1480));
   NOR2_X1 i_975 (.A1(n_1819), .A2(n_1807), .ZN(n_1481));
   NOR2_X1 i_976 (.A1(n_1819), .A2(n_1806), .ZN(n_1482));
   NOR2_X1 i_977 (.A1(n_1819), .A2(n_1805), .ZN(n_1483));
   NOR2_X1 i_978 (.A1(n_1819), .A2(n_1804), .ZN(n_1484));
   NOR2_X1 i_979 (.A1(n_1819), .A2(n_1803), .ZN(n_1485));
   NOR2_X1 i_980 (.A1(n_1819), .A2(n_1802), .ZN(n_1486));
   NOR2_X1 i_981 (.A1(n_1819), .A2(n_1801), .ZN(n_1487));
   NOR2_X1 i_982 (.A1(n_1819), .A2(n_1800), .ZN(n_1488));
   NOR2_X1 i_983 (.A1(n_1819), .A2(n_1799), .ZN(n_1489));
   NOR2_X1 i_984 (.A1(n_1819), .A2(n_1798), .ZN(n_1490));
   NOR2_X1 i_985 (.A1(n_1819), .A2(n_1797), .ZN(n_1491));
   NOR2_X1 i_986 (.A1(n_1819), .A2(n_1796), .ZN(n_1492));
   NOR2_X1 i_987 (.A1(n_1819), .A2(n_1795), .ZN(n_1493));
   NOR2_X1 i_988 (.A1(n_1819), .A2(n_1794), .ZN(n_1494));
   NOR2_X1 i_989 (.A1(n_1818), .A2(n_1816), .ZN(n_1495));
   NOR2_X1 i_990 (.A1(n_1818), .A2(n_1815), .ZN(n_1496));
   NOR2_X1 i_991 (.A1(n_1818), .A2(n_1814), .ZN(n_1497));
   NOR2_X1 i_992 (.A1(n_1818), .A2(n_1813), .ZN(n_1498));
   NOR2_X1 i_993 (.A1(n_1818), .A2(n_1812), .ZN(n_1499));
   NOR2_X1 i_994 (.A1(n_1818), .A2(n_1811), .ZN(n_1500));
   NOR2_X1 i_995 (.A1(n_1818), .A2(n_1810), .ZN(n_1501));
   NOR2_X1 i_996 (.A1(n_1818), .A2(n_1809), .ZN(n_1502));
   NOR2_X1 i_997 (.A1(n_1818), .A2(n_1808), .ZN(n_1503));
   NOR2_X1 i_998 (.A1(n_1818), .A2(n_1807), .ZN(n_1504));
   NOR2_X1 i_999 (.A1(n_1818), .A2(n_1806), .ZN(n_1505));
   NOR2_X1 i_1000 (.A1(n_1818), .A2(n_1805), .ZN(n_1506));
   NOR2_X1 i_1001 (.A1(n_1818), .A2(n_1804), .ZN(n_1507));
   NOR2_X1 i_1002 (.A1(n_1818), .A2(n_1803), .ZN(n_1508));
   NOR2_X1 i_1003 (.A1(n_1818), .A2(n_1802), .ZN(n_1509));
   NOR2_X1 i_1004 (.A1(n_1818), .A2(n_1801), .ZN(n_1510));
   NOR2_X1 i_1005 (.A1(n_1818), .A2(n_1800), .ZN(n_1511));
   NOR2_X1 i_1006 (.A1(n_1818), .A2(n_1799), .ZN(n_1512));
   NOR2_X1 i_1007 (.A1(n_1818), .A2(n_1798), .ZN(n_1513));
   NOR2_X1 i_1008 (.A1(n_1818), .A2(n_1797), .ZN(n_1514));
   NOR2_X1 i_1009 (.A1(n_1818), .A2(n_1796), .ZN(n_1515));
   NOR2_X1 i_1010 (.A1(n_1817), .A2(n_1816), .ZN(n_1516));
   NOR2_X1 i_1011 (.A1(n_1817), .A2(n_1815), .ZN(n_1517));
   NOR2_X1 i_1012 (.A1(n_1817), .A2(n_1814), .ZN(n_1518));
   NOR2_X1 i_1013 (.A1(n_1817), .A2(n_1813), .ZN(n_1519));
   NOR2_X1 i_1014 (.A1(n_1817), .A2(n_1812), .ZN(n_1520));
   NOR2_X1 i_1015 (.A1(n_1817), .A2(n_1811), .ZN(n_1521));
   NOR2_X1 i_1016 (.A1(n_1817), .A2(n_1810), .ZN(n_1522));
   NOR2_X1 i_1017 (.A1(n_1817), .A2(n_1809), .ZN(n_1523));
   NOR2_X1 i_1018 (.A1(n_1817), .A2(n_1808), .ZN(n_1524));
   NOR2_X1 i_1019 (.A1(n_1817), .A2(n_1807), .ZN(n_1525));
   NOR2_X1 i_1020 (.A1(n_1817), .A2(n_1806), .ZN(n_1526));
   NOR2_X1 i_1021 (.A1(n_1817), .A2(n_1805), .ZN(n_1527));
   NOR2_X1 i_1022 (.A1(n_1817), .A2(n_1804), .ZN(n_1528));
   NOR2_X1 i_1023 (.A1(n_1817), .A2(n_1803), .ZN(n_1529));
   NOR2_X1 i_1024 (.A1(n_1817), .A2(n_1802), .ZN(n_1530));
   NOR2_X1 i_1025 (.A1(n_1817), .A2(n_1801), .ZN(n_1531));
   NOR2_X1 i_1026 (.A1(n_1817), .A2(n_1800), .ZN(n_1532));
   NOR2_X1 i_1027 (.A1(n_1817), .A2(n_1799), .ZN(n_1533));
   NOR2_X1 i_1028 (.A1(n_1817), .A2(n_1798), .ZN(n_1534));
   NOR2_X1 i_1029 (.A1(n_1817), .A2(n_1797), .ZN(n_1535));
   INV_X1 i_1030 (.A(n_1536), .ZN(o_mantissa[1]));
   OAI21_X1 i_1031 (.A(n_1784), .B1(n_1787), .B2(n_1786), .ZN(n_1536));
   XOR2_X1 i_1032 (.A(n_1784), .B(n_1537), .Z(o_mantissa[2]));
   OAI21_X1 i_1033 (.A(n_1783), .B1(n_0), .B2(n_1789), .ZN(n_1537));
   XNOR2_X1 i_1034 (.A(n_1782), .B(n_1538), .ZN(o_mantissa[3]));
   OAI21_X1 i_1035 (.A(n_1790), .B1(n_2), .B2(n_4), .ZN(n_1538));
   XOR2_X1 i_1036 (.A(n_1780), .B(n_1539), .Z(o_mantissa[4]));
   XOR2_X1 i_1037 (.A(n_6), .B(n_10), .Z(n_1539));
   XOR2_X1 i_1038 (.A(n_1779), .B(n_1546), .Z(o_mantissa[5]));
   XOR2_X1 i_1039 (.A(n_1545), .B(n_1542), .Z(o_mantissa[6]));
   XOR2_X1 i_1040 (.A(n_1543), .B(n_1540), .Z(o_mantissa[7]));
   NOR2_X1 i_1041 (.A1(n_1776), .A2(n_1767), .ZN(n_1540));
   XNOR2_X1 i_1042 (.A(n_1547), .B(n_1541), .ZN(o_mantissa[8]));
   OAI22_X1 i_1043 (.A1(n_38), .A2(n_40), .B1(n_1767), .B2(n_1543), .ZN(n_1541));
   AOI21_X1 i_1044 (.A(n_1777), .B1(n_26), .B2(n_28), .ZN(n_1542));
   AOI21_X1 i_1045 (.A(n_1777), .B1(n_1771), .B2(n_1544), .ZN(n_1543));
   INV_X1 i_1046 (.A(n_1545), .ZN(n_1544));
   AOI21_X1 i_1047 (.A(n_1774), .B1(n_1779), .B2(n_1772), .ZN(n_1545));
   OAI21_X1 i_1048 (.A(n_1772), .B1(n_16), .B2(n_18), .ZN(n_1546));
   NOR2_X1 i_1049 (.A1(n_1778), .A2(n_1769), .ZN(n_1547));
   XOR2_X1 i_1050 (.A(n_1765), .B(n_1554), .Z(o_mantissa[9]));
   XOR2_X1 i_1051 (.A(n_1553), .B(n_1550), .Z(o_mantissa[10]));
   XOR2_X1 i_1052 (.A(n_1551), .B(n_1548), .Z(o_mantissa[11]));
   NOR2_X1 i_1053 (.A1(n_1762), .A2(n_1753), .ZN(n_1548));
   XNOR2_X1 i_1054 (.A(n_1555), .B(n_1549), .ZN(o_mantissa[12]));
   OAI22_X1 i_1055 (.A1(n_106), .A2(n_108), .B1(n_1753), .B2(n_1551), .ZN(n_1549));
   AOI21_X1 i_1056 (.A(n_1763), .B1(n_86), .B2(n_88), .ZN(n_1550));
   AOI21_X1 i_1057 (.A(n_1763), .B1(n_1757), .B2(n_1552), .ZN(n_1551));
   INV_X1 i_1058 (.A(n_1553), .ZN(n_1552));
   AOI21_X1 i_1059 (.A(n_1760), .B1(n_1765), .B2(n_1758), .ZN(n_1553));
   OAI21_X1 i_1060 (.A(n_1758), .B1(n_68), .B2(n_70), .ZN(n_1554));
   NOR2_X1 i_1061 (.A1(n_1764), .A2(n_1755), .ZN(n_1555));
   XOR2_X1 i_1062 (.A(n_1751), .B(n_1562), .Z(o_mantissa[13]));
   XOR2_X1 i_1063 (.A(n_1561), .B(n_1558), .Z(o_mantissa[14]));
   XOR2_X1 i_1064 (.A(n_1559), .B(n_1556), .Z(o_mantissa[15]));
   NOR2_X1 i_1065 (.A1(n_1748), .A2(n_1739), .ZN(n_1556));
   XNOR2_X1 i_1066 (.A(n_1563), .B(n_1557), .ZN(o_mantissa[16]));
   OAI22_X1 i_1067 (.A1(n_206), .A2(n_208), .B1(n_1739), .B2(n_1559), .ZN(n_1557));
   AOI21_X1 i_1068 (.A(n_1749), .B1(n_178), .B2(n_180), .ZN(n_1558));
   AOI21_X1 i_1069 (.A(n_1749), .B1(n_1743), .B2(n_1560), .ZN(n_1559));
   INV_X1 i_1070 (.A(n_1561), .ZN(n_1560));
   AOI21_X1 i_1071 (.A(n_1746), .B1(n_1751), .B2(n_1744), .ZN(n_1561));
   OAI21_X1 i_1072 (.A(n_1744), .B1(n_152), .B2(n_154), .ZN(n_1562));
   NOR2_X1 i_1073 (.A1(n_1750), .A2(n_1741), .ZN(n_1563));
   XOR2_X1 i_1074 (.A(n_1737), .B(n_1570), .Z(o_mantissa[17]));
   XOR2_X1 i_1075 (.A(n_1569), .B(n_1566), .Z(o_mantissa[18]));
   XOR2_X1 i_1076 (.A(n_1567), .B(n_1564), .Z(o_mantissa[19]));
   NOR2_X1 i_1077 (.A1(n_1706), .A2(n_1696), .ZN(n_1564));
   XNOR2_X1 i_1078 (.A(n_1571), .B(n_1565), .ZN(o_mantissa[20]));
   OAI21_X1 i_1079 (.A(n_1705), .B1(n_1696), .B2(n_1567), .ZN(n_1565));
   NOR2_X1 i_1080 (.A1(n_1708), .A2(n_1698), .ZN(n_1566));
   INV_X1 i_1081 (.A(n_1568), .ZN(n_1567));
   OAI21_X1 i_1082 (.A(n_1707), .B1(n_1698), .B2(n_1569), .ZN(n_1568));
   AOI21_X1 i_1083 (.A(n_1703), .B1(n_1737), .B2(n_1700), .ZN(n_1569));
   OAI21_X1 i_1084 (.A(n_1700), .B1(n_268), .B2(n_270), .ZN(n_1570));
   AOI21_X1 i_1085 (.A(n_1710), .B1(n_376), .B2(n_378), .ZN(n_1571));
   XOR2_X1 i_1086 (.A(n_1599), .B(n_1578), .Z(o_mantissa[21]));
   XOR2_X1 i_1087 (.A(n_1577), .B(n_1574), .Z(o_mantissa[22]));
   XOR2_X1 i_1088 (.A(n_1575), .B(n_1572), .Z(o_mantissa[23]));
   NOR2_X1 i_1089 (.A1(n_1731), .A2(n_1689), .ZN(n_1572));
   XNOR2_X1 i_1090 (.A(n_1579), .B(n_1573), .ZN(o_mantissa[24]));
   OAI21_X1 i_1091 (.A(n_1730), .B1(n_1689), .B2(n_1575), .ZN(n_1573));
   NOR2_X1 i_1092 (.A1(n_1733), .A2(n_1691), .ZN(n_1574));
   INV_X1 i_1093 (.A(n_1576), .ZN(n_1575));
   OAI21_X1 i_1094 (.A(n_1732), .B1(n_1691), .B2(n_1577), .ZN(n_1576));
   AOI21_X1 i_1095 (.A(n_1736), .B1(n_1693), .B2(n_1599), .ZN(n_1577));
   OAI21_X1 i_1096 (.A(n_1693), .B1(n_379), .B2(n_418), .ZN(n_1578));
   AOI21_X1 i_1097 (.A(n_1735), .B1(n_505), .B2(n_548), .ZN(n_1579));
   XOR2_X1 i_1098 (.A(n_1597), .B(n_1586), .Z(o_mantissa[25]));
   XOR2_X1 i_1099 (.A(n_1585), .B(n_1582), .Z(o_mantissa[26]));
   XOR2_X1 i_1100 (.A(n_1583), .B(n_1580), .Z(o_mantissa[27]));
   NOR2_X1 i_1101 (.A1(n_1717), .A2(n_1675), .ZN(n_1580));
   XNOR2_X1 i_1102 (.A(n_1587), .B(n_1581), .ZN(o_mantissa[28]));
   OAI21_X1 i_1103 (.A(n_1716), .B1(n_1675), .B2(n_1583), .ZN(n_1581));
   NOR2_X1 i_1104 (.A1(n_1719), .A2(n_1677), .ZN(n_1582));
   INV_X1 i_1105 (.A(n_1584), .ZN(n_1583));
   OAI21_X1 i_1106 (.A(n_1718), .B1(n_1677), .B2(n_1585), .ZN(n_1584));
   AOI21_X1 i_1107 (.A(n_1714), .B1(n_1679), .B2(n_1597), .ZN(n_1585));
   OAI21_X1 i_1108 (.A(n_1679), .B1(n_549), .B2(n_590), .ZN(n_1586));
   AOI21_X1 i_1109 (.A(n_1721), .B1(n_669), .B2(n_704), .ZN(n_1587));
   XNOR2_X1 i_1110 (.A(n_1596), .B(n_1595), .ZN(o_mantissa[29]));
   XOR2_X1 i_1111 (.A(n_1593), .B(n_1592), .Z(o_mantissa[30]));
   XNOR2_X1 i_1112 (.A(n_1589), .B(n_1588), .ZN(o_mantissa[31]));
   OAI22_X1 i_1113 (.A1(n_739), .A2(n_770), .B1(n_1685), .B2(n_1593), .ZN(n_1588));
   NOR2_X1 i_1114 (.A1(n_1725), .A2(n_1682), .ZN(n_1589));
   XNOR2_X1 i_1115 (.A(n_1601), .B(n_1590), .ZN(o_mantissa[32]));
   OAI21_X1 i_1116 (.A(n_1591), .B1(n_1724), .B2(n_1682), .ZN(n_1590));
   NAND3_X1 i_1117 (.A1(n_1683), .A2(n_1592), .A3(n_1594), .ZN(n_1591));
   NOR2_X1 i_1118 (.A1(n_1726), .A2(n_1685), .ZN(n_1592));
   INV_X1 i_1119 (.A(n_1594), .ZN(n_1593));
   OAI22_X1 i_1120 (.A1(n_705), .A2(n_738), .B1(n_1686), .B2(n_1596), .ZN(n_1594));
   OAI21_X1 i_1121 (.A(n_1687), .B1(n_705), .B2(n_738), .ZN(n_1595));
   OAI21_X1 i_1122 (.A(n_1674), .B1(n_1713), .B2(n_1597), .ZN(n_1596));
   INV_X1 i_1123 (.A(n_1598), .ZN(n_1597));
   OAI21_X1 i_1124 (.A(n_1688), .B1(n_1728), .B2(n_1599), .ZN(n_1598));
   INV_X1 i_1125 (.A(n_1600), .ZN(n_1599));
   OAI21_X1 i_1126 (.A(n_1695), .B1(n_1737), .B2(n_1702), .ZN(n_1600));
   AOI21_X1 i_1127 (.A(n_1727), .B1(n_801), .B2(n_828), .ZN(n_1601));
   XOR2_X1 i_1128 (.A(n_1672), .B(n_1608), .Z(o_mantissa[33]));
   XOR2_X1 i_1129 (.A(n_1607), .B(n_1604), .Z(o_mantissa[34]));
   XOR2_X1 i_1130 (.A(n_1605), .B(n_1602), .Z(o_mantissa[35]));
   NOR2_X1 i_1131 (.A1(n_1669), .A2(n_1660), .ZN(n_1602));
   XNOR2_X1 i_1132 (.A(n_1609), .B(n_1603), .ZN(o_mantissa[36]));
   OAI22_X1 i_1133 (.A1(n_879), .A2(n_900), .B1(n_1660), .B2(n_1605), .ZN(n_1603));
   AOI21_X1 i_1134 (.A(n_1670), .B1(n_855), .B2(n_878), .ZN(n_1604));
   AOI21_X1 i_1135 (.A(n_1670), .B1(n_1664), .B2(n_1606), .ZN(n_1605));
   INV_X1 i_1136 (.A(n_1607), .ZN(n_1606));
   AOI21_X1 i_1137 (.A(n_1667), .B1(n_1672), .B2(n_1665), .ZN(n_1607));
   OAI21_X1 i_1138 (.A(n_1665), .B1(n_829), .B2(n_854), .ZN(n_1608));
   NOR2_X1 i_1139 (.A1(n_1671), .A2(n_1662), .ZN(n_1609));
   XOR2_X1 i_1140 (.A(n_1658), .B(n_1616), .Z(o_mantissa[37]));
   XOR2_X1 i_1141 (.A(n_1615), .B(n_1612), .Z(o_mantissa[38]));
   XOR2_X1 i_1142 (.A(n_1613), .B(n_1610), .Z(o_mantissa[39]));
   NOR2_X1 i_1143 (.A1(n_1655), .A2(n_1646), .ZN(n_1610));
   XNOR2_X1 i_1144 (.A(n_1617), .B(n_1611), .ZN(o_mantissa[40]));
   OAI22_X1 i_1145 (.A1(n_955), .A2(n_968), .B1(n_1646), .B2(n_1613), .ZN(n_1611));
   AOI21_X1 i_1146 (.A(n_1656), .B1(n_939), .B2(n_954), .ZN(n_1612));
   AOI21_X1 i_1147 (.A(n_1656), .B1(n_1650), .B2(n_1614), .ZN(n_1613));
   INV_X1 i_1148 (.A(n_1615), .ZN(n_1614));
   AOI21_X1 i_1149 (.A(n_1653), .B1(n_1658), .B2(n_1651), .ZN(n_1615));
   OAI21_X1 i_1150 (.A(n_1651), .B1(n_921), .B2(n_938), .ZN(n_1616));
   NOR2_X1 i_1151 (.A1(n_1657), .A2(n_1648), .ZN(n_1617));
   XOR2_X1 i_1152 (.A(n_1644), .B(n_1624), .Z(o_mantissa[41]));
   XOR2_X1 i_1153 (.A(n_1623), .B(n_1622), .Z(o_mantissa[42]));
   XNOR2_X1 i_1154 (.A(n_1619), .B(n_1618), .ZN(o_mantissa[43]));
   OAI22_X1 i_1155 (.A1(n_991), .A2(n_998), .B1(n_1634), .B2(n_1623), .ZN(n_1618));
   NOR2_X1 i_1156 (.A1(n_1641), .A2(n_1630), .ZN(n_1619));
   XNOR2_X1 i_1157 (.A(n_1625), .B(n_1620), .ZN(o_mantissa[44]));
   OAI22_X1 i_1158 (.A1(n_1623), .A2(n_1621), .B1(n_1640), .B2(n_1630), .ZN(
      n_1620));
   NAND2_X1 i_1159 (.A1(n_1631), .A2(n_1622), .ZN(n_1621));
   NOR2_X1 i_1160 (.A1(n_1642), .A2(n_1634), .ZN(n_1622));
   AOI21_X1 i_1161 (.A(n_1638), .B1(n_1644), .B2(n_1636), .ZN(n_1623));
   OAI21_X1 i_1162 (.A(n_1636), .B1(n_981), .B2(n_990), .ZN(n_1624));
   NOR2_X1 i_1163 (.A1(n_1643), .A2(n_1632), .ZN(n_1625));
   XNOR2_X1 i_1164 (.A(n_1628), .B(n_1626), .ZN(o_mantissa[45]));
   AOI21_X1 i_1165 (.A(n_1792), .B1(n_1009), .B2(n_1010), .ZN(n_1626));
   XNOR2_X1 i_1166 (.A(n_1011), .B(n_1627), .ZN(o_mantissa[46]));
   OR2_X1 i_1167 (.A1(n_1011), .A2(n_1627), .ZN(o_mantissa[47]));
   OAI21_X1 i_1168 (.A(n_1793), .B1(n_1792), .B2(n_1628), .ZN(n_1627));
   NOR4_X1 i_1169 (.A1(n_1632), .A2(n_1629), .A3(n_1633), .A4(n_1637), .ZN(
      n_1628));
   NOR2_X1 i_1170 (.A1(n_1643), .A2(n_1631), .ZN(n_1629));
   INV_X1 i_1171 (.A(n_1631), .ZN(n_1630));
   NAND2_X1 i_1172 (.A1(n_999), .A2(n_1004), .ZN(n_1631));
   AND2_X1 i_1173 (.A1(n_1005), .A2(n_1008), .ZN(n_1632));
   AOI21_X1 i_1174 (.A(n_1639), .B1(n_1636), .B2(n_1635), .ZN(n_1633));
   INV_X1 i_1175 (.A(n_1635), .ZN(n_1634));
   NAND2_X1 i_1176 (.A1(n_991), .A2(n_998), .ZN(n_1635));
   NAND2_X1 i_1177 (.A1(n_981), .A2(n_990), .ZN(n_1636));
   NOR3_X1 i_1178 (.A1(n_1639), .A2(n_1638), .A3(n_1644), .ZN(n_1637));
   NOR2_X1 i_1179 (.A1(n_981), .A2(n_990), .ZN(n_1638));
   OAI21_X1 i_1180 (.A(n_1640), .B1(n_1005), .B2(n_1008), .ZN(n_1639));
   NOR2_X1 i_1181 (.A1(n_1642), .A2(n_1641), .ZN(n_1640));
   NOR2_X1 i_1182 (.A1(n_999), .A2(n_1004), .ZN(n_1641));
   NOR2_X1 i_1183 (.A1(n_991), .A2(n_998), .ZN(n_1642));
   NOR2_X1 i_1184 (.A1(n_1005), .A2(n_1008), .ZN(n_1643));
   NOR4_X1 i_1185 (.A1(n_1648), .A2(n_1645), .A3(n_1649), .A4(n_1652), .ZN(
      n_1644));
   NOR2_X1 i_1186 (.A1(n_1657), .A2(n_1647), .ZN(n_1645));
   INV_X1 i_1187 (.A(n_1647), .ZN(n_1646));
   NAND2_X1 i_1188 (.A1(n_955), .A2(n_968), .ZN(n_1647));
   AND2_X1 i_1189 (.A1(n_969), .A2(n_980), .ZN(n_1648));
   AOI21_X1 i_1190 (.A(n_1654), .B1(n_1651), .B2(n_1650), .ZN(n_1649));
   NAND2_X1 i_1191 (.A1(n_939), .A2(n_954), .ZN(n_1650));
   NAND2_X1 i_1192 (.A1(n_921), .A2(n_938), .ZN(n_1651));
   NOR3_X1 i_1193 (.A1(n_1654), .A2(n_1653), .A3(n_1658), .ZN(n_1652));
   NOR2_X1 i_1194 (.A1(n_921), .A2(n_938), .ZN(n_1653));
   OR3_X1 i_1195 (.A1(n_1657), .A2(n_1655), .A3(n_1656), .ZN(n_1654));
   NOR2_X1 i_1196 (.A1(n_955), .A2(n_968), .ZN(n_1655));
   NOR2_X1 i_1197 (.A1(n_939), .A2(n_954), .ZN(n_1656));
   NOR2_X1 i_1198 (.A1(n_969), .A2(n_980), .ZN(n_1657));
   NOR4_X1 i_1199 (.A1(n_1662), .A2(n_1659), .A3(n_1663), .A4(n_1666), .ZN(
      n_1658));
   NOR2_X1 i_1200 (.A1(n_1671), .A2(n_1661), .ZN(n_1659));
   INV_X1 i_1201 (.A(n_1661), .ZN(n_1660));
   NAND2_X1 i_1202 (.A1(n_879), .A2(n_900), .ZN(n_1661));
   AND2_X1 i_1203 (.A1(n_901), .A2(n_920), .ZN(n_1662));
   AOI21_X1 i_1204 (.A(n_1668), .B1(n_1665), .B2(n_1664), .ZN(n_1663));
   NAND2_X1 i_1205 (.A1(n_855), .A2(n_878), .ZN(n_1664));
   NAND2_X1 i_1206 (.A1(n_829), .A2(n_854), .ZN(n_1665));
   NOR3_X1 i_1207 (.A1(n_1668), .A2(n_1667), .A3(n_1672), .ZN(n_1666));
   NOR2_X1 i_1208 (.A1(n_829), .A2(n_854), .ZN(n_1667));
   OR3_X1 i_1209 (.A1(n_1671), .A2(n_1669), .A3(n_1670), .ZN(n_1668));
   NOR2_X1 i_1210 (.A1(n_879), .A2(n_900), .ZN(n_1669));
   NOR2_X1 i_1211 (.A1(n_855), .A2(n_878), .ZN(n_1670));
   NOR2_X1 i_1212 (.A1(n_901), .A2(n_920), .ZN(n_1671));
   NOR3_X1 i_1213 (.A1(n_1694), .A2(n_1673), .A3(n_1701), .ZN(n_1672));
   OAI221_X1 i_1214 (.A(n_1680), .B1(n_1722), .B2(n_1674), .C1(n_1712), .C2(
      n_1688), .ZN(n_1673));
   AOI221_X1 i_1215 (.A(n_1676), .B1(n_669), .B2(n_704), .C1(n_1720), .C2(n_1675), 
      .ZN(n_1674));
   AND2_X1 i_1216 (.A1(n_631), .A2(n_668), .ZN(n_1675));
   AOI21_X1 i_1217 (.A(n_1715), .B1(n_1679), .B2(n_1678), .ZN(n_1676));
   INV_X1 i_1218 (.A(n_1678), .ZN(n_1677));
   NAND2_X1 i_1219 (.A1(n_591), .A2(n_630), .ZN(n_1678));
   NAND2_X1 i_1220 (.A1(n_549), .A2(n_590), .ZN(n_1679));
   AOI21_X1 i_1221 (.A(n_1681), .B1(n_801), .B2(n_828), .ZN(n_1680));
   OAI21_X1 i_1222 (.A(n_1684), .B1(n_1727), .B2(n_1683), .ZN(n_1681));
   INV_X1 i_1223 (.A(n_1683), .ZN(n_1682));
   NAND2_X1 i_1224 (.A1(n_771), .A2(n_800), .ZN(n_1683));
   OAI21_X1 i_1225 (.A(n_1723), .B1(n_1686), .B2(n_1685), .ZN(n_1684));
   AND2_X1 i_1226 (.A1(n_739), .A2(n_770), .ZN(n_1685));
   INV_X1 i_1227 (.A(n_1687), .ZN(n_1686));
   NAND2_X1 i_1228 (.A1(n_705), .A2(n_738), .ZN(n_1687));
   AOI221_X1 i_1229 (.A(n_1690), .B1(n_505), .B2(n_548), .C1(n_1734), .C2(n_1689), 
      .ZN(n_1688));
   AND2_X1 i_1230 (.A1(n_461), .A2(n_504), .ZN(n_1689));
   AOI21_X1 i_1231 (.A(n_1729), .B1(n_1693), .B2(n_1692), .ZN(n_1690));
   INV_X1 i_1232 (.A(n_1692), .ZN(n_1691));
   NAND2_X1 i_1233 (.A1(n_419), .A2(n_460), .ZN(n_1692));
   NAND2_X1 i_1234 (.A1(n_379), .A2(n_418), .ZN(n_1693));
   NOR2_X1 i_1235 (.A1(n_1711), .A2(n_1695), .ZN(n_1694));
   AOI221_X1 i_1236 (.A(n_1697), .B1(n_376), .B2(n_378), .C1(n_1709), .C2(n_1696), 
      .ZN(n_1695));
   AND2_X1 i_1237 (.A1(n_305), .A2(n_340), .ZN(n_1696));
   AOI21_X1 i_1238 (.A(n_1704), .B1(n_1700), .B2(n_1699), .ZN(n_1697));
   INV_X1 i_1239 (.A(n_1699), .ZN(n_1698));
   NAND2_X1 i_1240 (.A1(n_271), .A2(n_304), .ZN(n_1699));
   NAND2_X1 i_1241 (.A1(n_268), .A2(n_270), .ZN(n_1700));
   NOR3_X1 i_1242 (.A1(n_1711), .A2(n_1702), .A3(n_1737), .ZN(n_1701));
   OR2_X1 i_1243 (.A1(n_1704), .A2(n_1703), .ZN(n_1702));
   NOR2_X1 i_1244 (.A1(n_268), .A2(n_270), .ZN(n_1703));
   NAND3_X1 i_1245 (.A1(n_1709), .A2(n_1705), .A3(n_1707), .ZN(n_1704));
   INV_X1 i_1246 (.A(n_1706), .ZN(n_1705));
   NOR2_X1 i_1247 (.A1(n_305), .A2(n_340), .ZN(n_1706));
   INV_X1 i_1248 (.A(n_1708), .ZN(n_1707));
   NOR2_X1 i_1249 (.A1(n_271), .A2(n_304), .ZN(n_1708));
   INV_X1 i_1250 (.A(n_1710), .ZN(n_1709));
   NOR2_X1 i_1251 (.A1(n_376), .A2(n_378), .ZN(n_1710));
   OR2_X1 i_1252 (.A1(n_1728), .A2(n_1712), .ZN(n_1711));
   OR2_X1 i_1253 (.A1(n_1722), .A2(n_1713), .ZN(n_1712));
   OR2_X1 i_1254 (.A1(n_1715), .A2(n_1714), .ZN(n_1713));
   NOR2_X1 i_1255 (.A1(n_549), .A2(n_590), .ZN(n_1714));
   NAND3_X1 i_1256 (.A1(n_1720), .A2(n_1716), .A3(n_1718), .ZN(n_1715));
   INV_X1 i_1257 (.A(n_1717), .ZN(n_1716));
   NOR2_X1 i_1258 (.A1(n_631), .A2(n_668), .ZN(n_1717));
   INV_X1 i_1259 (.A(n_1719), .ZN(n_1718));
   NOR2_X1 i_1260 (.A1(n_591), .A2(n_630), .ZN(n_1719));
   INV_X1 i_1261 (.A(n_1721), .ZN(n_1720));
   NOR2_X1 i_1262 (.A1(n_669), .A2(n_704), .ZN(n_1721));
   OAI21_X1 i_1263 (.A(n_1723), .B1(n_705), .B2(n_738), .ZN(n_1722));
   NOR3_X1 i_1264 (.A1(n_1727), .A2(n_1725), .A3(n_1726), .ZN(n_1723));
   NOR2_X1 i_1265 (.A1(n_1726), .A2(n_1725), .ZN(n_1724));
   NOR2_X1 i_1266 (.A1(n_771), .A2(n_800), .ZN(n_1725));
   NOR2_X1 i_1267 (.A1(n_739), .A2(n_770), .ZN(n_1726));
   NOR2_X1 i_1268 (.A1(n_801), .A2(n_828), .ZN(n_1727));
   OR2_X1 i_1269 (.A1(n_1736), .A2(n_1729), .ZN(n_1728));
   NAND3_X1 i_1270 (.A1(n_1734), .A2(n_1730), .A3(n_1732), .ZN(n_1729));
   INV_X1 i_1271 (.A(n_1731), .ZN(n_1730));
   NOR2_X1 i_1272 (.A1(n_461), .A2(n_504), .ZN(n_1731));
   INV_X1 i_1273 (.A(n_1733), .ZN(n_1732));
   NOR2_X1 i_1274 (.A1(n_419), .A2(n_460), .ZN(n_1733));
   INV_X1 i_1275 (.A(n_1735), .ZN(n_1734));
   NOR2_X1 i_1276 (.A1(n_505), .A2(n_548), .ZN(n_1735));
   NOR2_X1 i_1277 (.A1(n_379), .A2(n_418), .ZN(n_1736));
   NOR4_X1 i_1278 (.A1(n_1741), .A2(n_1738), .A3(n_1742), .A4(n_1745), .ZN(
      n_1737));
   NOR2_X1 i_1279 (.A1(n_1750), .A2(n_1740), .ZN(n_1738));
   INV_X1 i_1280 (.A(n_1740), .ZN(n_1739));
   NAND2_X1 i_1281 (.A1(n_206), .A2(n_208), .ZN(n_1740));
   AND2_X1 i_1282 (.A1(n_236), .A2(n_238), .ZN(n_1741));
   AOI21_X1 i_1283 (.A(n_1747), .B1(n_1744), .B2(n_1743), .ZN(n_1742));
   NAND2_X1 i_1284 (.A1(n_178), .A2(n_180), .ZN(n_1743));
   NAND2_X1 i_1285 (.A1(n_152), .A2(n_154), .ZN(n_1744));
   NOR3_X1 i_1286 (.A1(n_1747), .A2(n_1746), .A3(n_1751), .ZN(n_1745));
   NOR2_X1 i_1287 (.A1(n_152), .A2(n_154), .ZN(n_1746));
   OR3_X1 i_1288 (.A1(n_1750), .A2(n_1748), .A3(n_1749), .ZN(n_1747));
   NOR2_X1 i_1289 (.A1(n_206), .A2(n_208), .ZN(n_1748));
   NOR2_X1 i_1290 (.A1(n_178), .A2(n_180), .ZN(n_1749));
   NOR2_X1 i_1291 (.A1(n_236), .A2(n_238), .ZN(n_1750));
   NOR4_X1 i_1292 (.A1(n_1755), .A2(n_1752), .A3(n_1756), .A4(n_1759), .ZN(
      n_1751));
   NOR2_X1 i_1293 (.A1(n_1764), .A2(n_1754), .ZN(n_1752));
   INV_X1 i_1294 (.A(n_1754), .ZN(n_1753));
   NAND2_X1 i_1295 (.A1(n_106), .A2(n_108), .ZN(n_1754));
   AND2_X1 i_1296 (.A1(n_128), .A2(n_130), .ZN(n_1755));
   AOI21_X1 i_1297 (.A(n_1761), .B1(n_1758), .B2(n_1757), .ZN(n_1756));
   NAND2_X1 i_1298 (.A1(n_86), .A2(n_88), .ZN(n_1757));
   NAND2_X1 i_1299 (.A1(n_68), .A2(n_70), .ZN(n_1758));
   NOR3_X1 i_1300 (.A1(n_1761), .A2(n_1760), .A3(n_1765), .ZN(n_1759));
   NOR2_X1 i_1301 (.A1(n_68), .A2(n_70), .ZN(n_1760));
   OR3_X1 i_1302 (.A1(n_1764), .A2(n_1762), .A3(n_1763), .ZN(n_1761));
   NOR2_X1 i_1303 (.A1(n_106), .A2(n_108), .ZN(n_1762));
   NOR2_X1 i_1304 (.A1(n_86), .A2(n_88), .ZN(n_1763));
   NOR2_X1 i_1305 (.A1(n_128), .A2(n_130), .ZN(n_1764));
   NOR4_X1 i_1306 (.A1(n_1769), .A2(n_1766), .A3(n_1770), .A4(n_1773), .ZN(
      n_1765));
   NOR2_X1 i_1307 (.A1(n_1778), .A2(n_1768), .ZN(n_1766));
   INV_X1 i_1308 (.A(n_1768), .ZN(n_1767));
   NAND2_X1 i_1309 (.A1(n_38), .A2(n_40), .ZN(n_1768));
   AND2_X1 i_1310 (.A1(n_52), .A2(n_54), .ZN(n_1769));
   AOI21_X1 i_1311 (.A(n_1775), .B1(n_1772), .B2(n_1771), .ZN(n_1770));
   NAND2_X1 i_1312 (.A1(n_26), .A2(n_28), .ZN(n_1771));
   NAND2_X1 i_1313 (.A1(n_16), .A2(n_18), .ZN(n_1772));
   NOR3_X1 i_1314 (.A1(n_1775), .A2(n_1774), .A3(n_1779), .ZN(n_1773));
   NOR2_X1 i_1315 (.A1(n_16), .A2(n_18), .ZN(n_1774));
   OR3_X1 i_1316 (.A1(n_1778), .A2(n_1776), .A3(n_1777), .ZN(n_1775));
   NOR2_X1 i_1317 (.A1(n_38), .A2(n_40), .ZN(n_1776));
   NOR2_X1 i_1318 (.A1(n_26), .A2(n_28), .ZN(n_1777));
   NOR2_X1 i_1319 (.A1(n_52), .A2(n_54), .ZN(n_1778));
   OAI22_X1 i_1320 (.A1(n_6), .A2(n_10), .B1(n_1791), .B2(n_1780), .ZN(n_1779));
   NAND2_X1 i_1321 (.A1(n_1790), .A2(n_1781), .ZN(n_1780));
   OAI21_X1 i_1322 (.A(n_1782), .B1(n_2), .B2(n_4), .ZN(n_1781));
   AOI21_X1 i_1323 (.A(n_1788), .B1(n_1784), .B2(n_1783), .ZN(n_1782));
   NAND2_X1 i_1324 (.A1(n_0), .A2(n_1789), .ZN(n_1783));
   NAND2_X1 i_1325 (.A1(o_mantissa[0]), .A2(n_1785), .ZN(n_1784));
   NOR2_X1 i_1326 (.A1(n_1818), .A2(n_1795), .ZN(n_1785));
   NOR2_X1 i_1327 (.A1(n_1817), .A2(n_1794), .ZN(o_mantissa[0]));
   NOR2_X1 i_1328 (.A1(n_1817), .A2(n_1795), .ZN(n_1786));
   NOR2_X1 i_1329 (.A1(n_1818), .A2(n_1794), .ZN(n_1787));
   NOR2_X1 i_1330 (.A1(n_0), .A2(n_1789), .ZN(n_1788));
   NOR2_X1 i_1331 (.A1(n_1817), .A2(n_1796), .ZN(n_1789));
   NAND2_X1 i_1332 (.A1(n_2), .A2(n_4), .ZN(n_1790));
   AND2_X1 i_1333 (.A1(n_6), .A2(n_10), .ZN(n_1791));
   NOR2_X1 i_1334 (.A1(n_1009), .A2(n_1010), .ZN(n_1792));
   NAND2_X1 i_1335 (.A1(n_1009), .A2(n_1010), .ZN(n_1793));
   INV_X1 i_1336 (.A(a_mantissa[0]), .ZN(n_1794));
   INV_X1 i_1337 (.A(a_mantissa[1]), .ZN(n_1795));
   INV_X1 i_1338 (.A(a_mantissa[2]), .ZN(n_1796));
   INV_X1 i_1339 (.A(a_mantissa[3]), .ZN(n_1797));
   INV_X1 i_1340 (.A(a_mantissa[4]), .ZN(n_1798));
   INV_X1 i_1341 (.A(a_mantissa[5]), .ZN(n_1799));
   INV_X1 i_1342 (.A(a_mantissa[6]), .ZN(n_1800));
   INV_X1 i_1343 (.A(a_mantissa[7]), .ZN(n_1801));
   INV_X1 i_1344 (.A(a_mantissa[8]), .ZN(n_1802));
   INV_X1 i_1345 (.A(a_mantissa[9]), .ZN(n_1803));
   INV_X1 i_1346 (.A(a_mantissa[10]), .ZN(n_1804));
   INV_X1 i_1347 (.A(a_mantissa[11]), .ZN(n_1805));
   INV_X1 i_1348 (.A(a_mantissa[12]), .ZN(n_1806));
   INV_X1 i_1349 (.A(a_mantissa[13]), .ZN(n_1807));
   INV_X1 i_1350 (.A(a_mantissa[14]), .ZN(n_1808));
   INV_X1 i_1351 (.A(a_mantissa[15]), .ZN(n_1809));
   INV_X1 i_1352 (.A(a_mantissa[16]), .ZN(n_1810));
   INV_X1 i_1353 (.A(a_mantissa[17]), .ZN(n_1811));
   INV_X1 i_1354 (.A(a_mantissa[18]), .ZN(n_1812));
   INV_X1 i_1355 (.A(a_mantissa[19]), .ZN(n_1813));
   INV_X1 i_1356 (.A(a_mantissa[20]), .ZN(n_1814));
   INV_X1 i_1357 (.A(a_mantissa[21]), .ZN(n_1815));
   INV_X1 i_1358 (.A(a_mantissa[22]), .ZN(n_1816));
   INV_X1 i_1359 (.A(b_mantissa[0]), .ZN(n_1817));
   INV_X1 i_1360 (.A(b_mantissa[1]), .ZN(n_1818));
   INV_X1 i_1361 (.A(b_mantissa[2]), .ZN(n_1819));
   INV_X1 i_1362 (.A(b_mantissa[3]), .ZN(n_1820));
   INV_X1 i_1363 (.A(b_mantissa[4]), .ZN(n_1821));
   INV_X1 i_1364 (.A(b_mantissa[5]), .ZN(n_1822));
   INV_X1 i_1365 (.A(b_mantissa[6]), .ZN(n_1823));
   INV_X1 i_1366 (.A(b_mantissa[7]), .ZN(n_1824));
   INV_X1 i_1367 (.A(b_mantissa[8]), .ZN(n_1825));
   INV_X1 i_1368 (.A(b_mantissa[9]), .ZN(n_1826));
   INV_X1 i_1369 (.A(b_mantissa[10]), .ZN(n_1827));
   INV_X1 i_1370 (.A(b_mantissa[11]), .ZN(n_1828));
   INV_X1 i_1371 (.A(b_mantissa[12]), .ZN(n_1829));
   INV_X1 i_1372 (.A(b_mantissa[13]), .ZN(n_1830));
   INV_X1 i_1373 (.A(b_mantissa[14]), .ZN(n_1831));
   INV_X1 i_1374 (.A(b_mantissa[15]), .ZN(n_1832));
   INV_X1 i_1375 (.A(b_mantissa[16]), .ZN(n_1833));
   INV_X1 i_1376 (.A(b_mantissa[17]), .ZN(n_1834));
   INV_X1 i_1377 (.A(b_mantissa[18]), .ZN(n_1835));
   INV_X1 i_1378 (.A(b_mantissa[19]), .ZN(n_1836));
   INV_X1 i_1379 (.A(b_mantissa[20]), .ZN(n_1837));
   INV_X1 i_1380 (.A(b_mantissa[21]), .ZN(n_1838));
   INV_X1 i_1381 (.A(b_mantissa[22]), .ZN(n_1839));
endmodule

module datapath__0_5(p_0, p_1, O_final_mantessa);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]O_final_mantessa;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(O_final_mantessa[0]));
   HA_X1 i_1 (.A(p_1[1]), .B(n_0), .CO(n_1), .S(O_final_mantessa[1]));
   HA_X1 i_2 (.A(p_1[2]), .B(n_1), .CO(n_2), .S(O_final_mantessa[2]));
   HA_X1 i_3 (.A(p_1[3]), .B(n_2), .CO(n_3), .S(O_final_mantessa[3]));
   HA_X1 i_4 (.A(p_1[4]), .B(n_3), .CO(n_4), .S(O_final_mantessa[4]));
   HA_X1 i_5 (.A(p_1[5]), .B(n_4), .CO(n_5), .S(O_final_mantessa[5]));
   HA_X1 i_6 (.A(p_1[6]), .B(n_5), .CO(n_6), .S(O_final_mantessa[6]));
   HA_X1 i_7 (.A(p_1[7]), .B(n_6), .CO(n_7), .S(O_final_mantessa[7]));
   HA_X1 i_8 (.A(p_1[8]), .B(n_7), .CO(n_8), .S(O_final_mantessa[8]));
   HA_X1 i_9 (.A(p_1[9]), .B(n_8), .CO(n_9), .S(O_final_mantessa[9]));
   HA_X1 i_10 (.A(p_1[10]), .B(n_9), .CO(n_10), .S(O_final_mantessa[10]));
   HA_X1 i_11 (.A(p_1[11]), .B(n_10), .CO(n_11), .S(O_final_mantessa[11]));
   HA_X1 i_12 (.A(p_1[12]), .B(n_11), .CO(n_12), .S(O_final_mantessa[12]));
   HA_X1 i_13 (.A(p_1[13]), .B(n_12), .CO(n_13), .S(O_final_mantessa[13]));
   HA_X1 i_14 (.A(p_1[14]), .B(n_13), .CO(n_14), .S(O_final_mantessa[14]));
   HA_X1 i_15 (.A(p_1[15]), .B(n_14), .CO(n_15), .S(O_final_mantessa[15]));
   HA_X1 i_16 (.A(p_1[16]), .B(n_15), .CO(n_16), .S(O_final_mantessa[16]));
   HA_X1 i_17 (.A(p_1[17]), .B(n_16), .CO(n_17), .S(O_final_mantessa[17]));
   HA_X1 i_18 (.A(p_1[18]), .B(n_17), .CO(n_18), .S(O_final_mantessa[18]));
   HA_X1 i_19 (.A(p_1[19]), .B(n_18), .CO(n_19), .S(O_final_mantessa[19]));
   HA_X1 i_20 (.A(p_1[20]), .B(n_19), .CO(n_20), .S(O_final_mantessa[20]));
   HA_X1 i_21 (.A(p_1[21]), .B(n_20), .CO(n_21), .S(O_final_mantessa[21]));
   XOR2_X1 i_22 (.A(p_1[22]), .B(n_21), .Z(O_final_mantessa[22]));
endmodule

module FloatingPointMultiplier(A, B, O, OF);
   input [31:0]A;
   input [31:0]B;
   output [31:0]O;
   output OF;

   wire [47:0]o_mantissa;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;
   wire n_1_10;
   wire n_1_11;
   wire n_1_12;
   wire n_1_13;
   wire n_1_15;
   wire n_1_16;
   wire n_1_24;
   wire n_1_17;
   wire n_1_25;
   wire n_1_18;
   wire n_1_26;
   wire n_1_19;
   wire n_1_27;
   wire n_1_20;
   wire n_1_28;
   wire n_1_21;
   wire n_1_29;
   wire n_1_22;
   wire n_1_30;
   wire n_1_23;
   wire n_1_14;
   wire n_1_0;
   wire n_1_1;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_53;
   wire n_1_54;
   wire n_1_55;
   wire n_1_56;
   wire n_1_57;
   wire n_1_58;
   wire n_1_59;
   wire n_1_60;
   wire n_1_61;
   wire n_1_62;
   wire n_1_63;
   wire n_1_64;
   wire n_1_74;
   wire n_1_75;
   wire n_1_76;
   wire n_1_77;
   wire n_1_78;
   wire n_1_79;
   wire n_1_80;
   wire n_1_81;
   wire n_1_82;
   wire n_1_83;
   wire n_1_84;
   wire n_1_85;
   wire n_1_86;
   wire n_1_87;
   wire n_1_88;
   wire n_1_89;
   wire n_1_90;
   wire n_1_91;
   wire n_1_92;
   wire n_1_93;
   wire n_1_94;
   wire n_1_95;
   wire n_1_96;
   wire n_1_97;
   wire n_1_98;
   wire n_1_99;
   wire n_1_100;
   wire n_1_101;
   wire n_1_102;
   wire n_1_103;
   wire n_1_104;
   wire n_1_65;
   wire n_1_66;
   wire n_1_67;
   wire n_1_68;
   wire n_1_69;
   wire n_1_70;
   wire n_1_71;
   wire n_1_72;
   wire n_1_73;
   wire n_1_105;

   datapath i_0 (.b_mantissa({uc_0, B[22], B[21], B[20], B[19], B[18], B[17], 
      B[16], B[15], B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], 
      B[5], B[4], B[3], B[2], B[1], B[0]}), .a_mantissa({uc_1, A[22], A[21], 
      A[20], A[19], A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], 
      A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0]}), 
      .o_mantissa(o_mantissa));
   datapath__0_5 i_5 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, n_46}), .p_1({n_45, n_44, n_43, n_42, n_41, n_40, n_39, n_38, n_37, 
      n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, n_28, n_27, n_26, n_25, 
      n_24, n_23}), .O_final_mantessa({n_22, n_21, n_20, n_19, n_18, n_17, n_16, 
      n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7, n_6, n_5, n_4, n_3, n_2, 
      n_1, n_0}));
   HA_X1 i_1_0 (.A(B[24]), .B(A[24]), .CO(n_1_3), .S(n_1_2));
   HA_X1 i_1_1 (.A(B[25]), .B(A[25]), .CO(n_1_5), .S(n_1_4));
   HA_X1 i_1_2 (.A(B[26]), .B(A[26]), .CO(n_1_7), .S(n_1_6));
   HA_X1 i_1_3 (.A(B[27]), .B(A[27]), .CO(n_1_9), .S(n_1_8));
   HA_X1 i_1_4 (.A(B[28]), .B(A[28]), .CO(n_1_11), .S(n_1_10));
   HA_X1 i_1_5 (.A(B[29]), .B(A[29]), .CO(n_1_13), .S(n_1_12));
   HA_X1 i_1_6 (.A(A[23]), .B(n_1_0), .CO(n_1_16), .S(n_1_15));
   FA_X1 i_1_7 (.A(n_1_1), .B(n_1_2), .CI(n_1_16), .CO(n_1_17), .S(n_1_24));
   FA_X1 i_1_8 (.A(n_1_3), .B(n_1_4), .CI(n_1_17), .CO(n_1_18), .S(n_1_25));
   FA_X1 i_1_9 (.A(n_1_5), .B(n_1_6), .CI(n_1_18), .CO(n_1_19), .S(n_1_26));
   FA_X1 i_1_10 (.A(n_1_7), .B(n_1_8), .CI(n_1_19), .CO(n_1_20), .S(n_1_27));
   FA_X1 i_1_11 (.A(n_1_9), .B(n_1_10), .CI(n_1_20), .CO(n_1_21), .S(n_1_28));
   FA_X1 i_1_12 (.A(n_1_11), .B(n_1_12), .CI(n_1_21), .CO(n_1_22), .S(n_1_29));
   FA_X1 i_1_13 (.A(n_1_13), .B(n_1_14), .CI(n_1_22), .CO(n_1_23), .S(n_1_30));
   XNOR2_X1 i_1_14 (.A(B[30]), .B(A[30]), .ZN(n_1_14));
   XNOR2_X1 i_1_15 (.A(B[23]), .B(o_mantissa[47]), .ZN(n_1_0));
   OR2_X1 i_1_16 (.A1(B[23]), .A2(o_mantissa[47]), .ZN(n_1_1));
   NOR2_X1 i_1_17 (.A1(n_1_33), .A2(n_1_31), .ZN(OF));
   XNOR2_X1 i_1_18 (.A(n_1_23), .B(n_1_32), .ZN(n_1_31));
   NOR2_X1 i_1_19 (.A1(B[30]), .A2(A[30]), .ZN(n_1_32));
   OAI21_X1 i_1_20 (.A(n_1_34), .B1(n_1_33), .B2(n_1_82), .ZN(O[0]));
   OAI21_X1 i_1_21 (.A(n_1_34), .B1(n_1_33), .B2(n_1_83), .ZN(O[1]));
   OAI21_X1 i_1_22 (.A(n_1_34), .B1(n_1_33), .B2(n_1_84), .ZN(O[2]));
   OAI21_X1 i_1_23 (.A(n_1_34), .B1(n_1_33), .B2(n_1_85), .ZN(O[3]));
   OAI21_X1 i_1_24 (.A(n_1_34), .B1(n_1_33), .B2(n_1_86), .ZN(O[4]));
   OAI21_X1 i_1_25 (.A(n_1_34), .B1(n_1_33), .B2(n_1_87), .ZN(O[5]));
   OAI21_X1 i_1_26 (.A(n_1_34), .B1(n_1_33), .B2(n_1_88), .ZN(O[6]));
   OAI21_X1 i_1_27 (.A(n_1_34), .B1(n_1_33), .B2(n_1_89), .ZN(O[7]));
   OAI21_X1 i_1_28 (.A(n_1_34), .B1(n_1_33), .B2(n_1_90), .ZN(O[8]));
   OAI21_X1 i_1_29 (.A(n_1_34), .B1(n_1_33), .B2(n_1_91), .ZN(O[9]));
   OAI21_X1 i_1_30 (.A(n_1_34), .B1(n_1_33), .B2(n_1_92), .ZN(O[10]));
   OAI21_X1 i_1_31 (.A(n_1_34), .B1(n_1_33), .B2(n_1_93), .ZN(O[11]));
   OAI21_X1 i_1_32 (.A(n_1_34), .B1(n_1_33), .B2(n_1_94), .ZN(O[12]));
   OAI21_X1 i_1_33 (.A(n_1_34), .B1(n_1_33), .B2(n_1_95), .ZN(O[13]));
   OAI21_X1 i_1_34 (.A(n_1_34), .B1(n_1_33), .B2(n_1_96), .ZN(O[14]));
   OAI21_X1 i_1_35 (.A(n_1_34), .B1(n_1_33), .B2(n_1_97), .ZN(O[15]));
   OAI21_X1 i_1_36 (.A(n_1_34), .B1(n_1_33), .B2(n_1_98), .ZN(O[16]));
   OAI21_X1 i_1_37 (.A(n_1_34), .B1(n_1_33), .B2(n_1_99), .ZN(O[17]));
   OAI21_X1 i_1_38 (.A(n_1_34), .B1(n_1_33), .B2(n_1_100), .ZN(O[18]));
   OAI21_X1 i_1_39 (.A(n_1_34), .B1(n_1_33), .B2(n_1_101), .ZN(O[19]));
   OAI21_X1 i_1_40 (.A(n_1_34), .B1(n_1_33), .B2(n_1_102), .ZN(O[20]));
   OAI21_X1 i_1_41 (.A(n_1_34), .B1(n_1_33), .B2(n_1_103), .ZN(O[21]));
   OAI21_X1 i_1_42 (.A(n_1_34), .B1(n_1_33), .B2(n_1_104), .ZN(O[22]));
   NAND2_X1 i_1_43 (.A1(n_1_58), .A2(n_1_36), .ZN(n_1_33));
   AOI221_X1 i_1_44 (.A(n_1_35), .B1(n_1_40), .B2(n_1_59), .C1(n_1_62), .C2(
      n_1_50), .ZN(n_1_34));
   NOR2_X1 i_1_45 (.A1(n_1_58), .A2(n_1_36), .ZN(n_1_35));
   OAI21_X1 i_1_46 (.A(n_1_58), .B1(n_1_37), .B2(n_1_81), .ZN(O[23]));
   OAI21_X1 i_1_47 (.A(n_1_58), .B1(n_1_37), .B2(n_1_80), .ZN(O[24]));
   OAI21_X1 i_1_48 (.A(n_1_58), .B1(n_1_37), .B2(n_1_79), .ZN(O[25]));
   OAI21_X1 i_1_49 (.A(n_1_58), .B1(n_1_37), .B2(n_1_78), .ZN(O[26]));
   OAI21_X1 i_1_50 (.A(n_1_58), .B1(n_1_37), .B2(n_1_77), .ZN(O[27]));
   OAI21_X1 i_1_51 (.A(n_1_58), .B1(n_1_37), .B2(n_1_76), .ZN(O[28]));
   OAI21_X1 i_1_52 (.A(n_1_58), .B1(n_1_37), .B2(n_1_75), .ZN(O[29]));
   OAI21_X1 i_1_53 (.A(n_1_58), .B1(n_1_37), .B2(n_1_74), .ZN(O[30]));
   INV_X1 i_1_54 (.A(n_1_37), .ZN(n_1_36));
   OAI33_X1 i_1_55 (.A1(n_1_50), .A2(n_1_49), .A3(n_1_48), .B1(n_1_40), .B2(
      n_1_39), .B3(n_1_38), .ZN(n_1_37));
   OR4_X1 i_1_56 (.A1(B[29]), .A2(B[28]), .A3(B[27]), .A4(B[26]), .ZN(n_1_38));
   OR4_X1 i_1_57 (.A1(B[30]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_1_39));
   NAND3_X1 i_1_58 (.A1(n_1_45), .A2(n_1_44), .A3(n_1_41), .ZN(n_1_40));
   AND4_X1 i_1_59 (.A1(n_1_47), .A2(n_1_46), .A3(n_1_43), .A4(n_1_42), .ZN(
      n_1_41));
   NOR4_X1 i_1_60 (.A1(B[6]), .A2(B[3]), .A3(B[2]), .A4(B[0]), .ZN(n_1_42));
   NOR4_X1 i_1_61 (.A1(B[13]), .A2(B[12]), .A3(B[10]), .A4(B[7]), .ZN(n_1_43));
   NOR3_X1 i_1_62 (.A1(B[5]), .A2(B[4]), .A3(B[1]), .ZN(n_1_44));
   NOR4_X1 i_1_63 (.A1(B[14]), .A2(B[11]), .A3(B[9]), .A4(B[8]), .ZN(n_1_45));
   NOR4_X1 i_1_64 (.A1(B[22]), .A2(B[19]), .A3(B[17]), .A4(B[16]), .ZN(n_1_46));
   NOR4_X1 i_1_65 (.A1(B[21]), .A2(B[20]), .A3(B[18]), .A4(B[15]), .ZN(n_1_47));
   OR4_X1 i_1_66 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_1_48));
   OR4_X1 i_1_67 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_1_49));
   NAND3_X1 i_1_68 (.A1(n_1_55), .A2(n_1_54), .A3(n_1_51), .ZN(n_1_50));
   AND4_X1 i_1_69 (.A1(n_1_57), .A2(n_1_56), .A3(n_1_53), .A4(n_1_52), .ZN(
      n_1_51));
   NOR4_X1 i_1_70 (.A1(A[6]), .A2(A[3]), .A3(A[2]), .A4(A[0]), .ZN(n_1_52));
   NOR4_X1 i_1_71 (.A1(A[13]), .A2(A[12]), .A3(A[10]), .A4(A[7]), .ZN(n_1_53));
   NOR3_X1 i_1_72 (.A1(A[5]), .A2(A[4]), .A3(A[1]), .ZN(n_1_54));
   NOR4_X1 i_1_73 (.A1(A[14]), .A2(A[11]), .A3(A[9]), .A4(A[8]), .ZN(n_1_55));
   NOR4_X1 i_1_74 (.A1(A[22]), .A2(A[19]), .A3(A[17]), .A4(A[16]), .ZN(n_1_56));
   NOR4_X1 i_1_75 (.A1(A[21]), .A2(A[20]), .A3(A[18]), .A4(A[15]), .ZN(n_1_57));
   NOR2_X1 i_1_76 (.A1(n_1_62), .A2(n_1_59), .ZN(n_1_58));
   NOR2_X1 i_1_77 (.A1(n_1_61), .A2(n_1_60), .ZN(n_1_59));
   NAND4_X1 i_1_78 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_1_60));
   NAND4_X1 i_1_79 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(n_1_61));
   NOR2_X1 i_1_80 (.A1(n_1_64), .A2(n_1_63), .ZN(n_1_62));
   NAND4_X1 i_1_81 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_1_63));
   NAND4_X1 i_1_82 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_1_64));
   XOR2_X1 i_1_83 (.A(B[31]), .B(A[31]), .Z(O[31]));
   MUX2_X1 i_1_94 (.A(o_mantissa[23]), .B(o_mantissa[24]), .S(o_mantissa[47]), 
      .Z(n_23));
   MUX2_X1 i_1_95 (.A(o_mantissa[24]), .B(o_mantissa[25]), .S(o_mantissa[47]), 
      .Z(n_24));
   MUX2_X1 i_1_96 (.A(o_mantissa[25]), .B(o_mantissa[26]), .S(o_mantissa[47]), 
      .Z(n_25));
   MUX2_X1 i_1_97 (.A(o_mantissa[26]), .B(o_mantissa[27]), .S(o_mantissa[47]), 
      .Z(n_26));
   MUX2_X1 i_1_98 (.A(o_mantissa[27]), .B(o_mantissa[28]), .S(o_mantissa[47]), 
      .Z(n_27));
   MUX2_X1 i_1_99 (.A(o_mantissa[28]), .B(o_mantissa[29]), .S(o_mantissa[47]), 
      .Z(n_28));
   MUX2_X1 i_1_100 (.A(o_mantissa[29]), .B(o_mantissa[30]), .S(o_mantissa[47]), 
      .Z(n_29));
   MUX2_X1 i_1_101 (.A(o_mantissa[30]), .B(o_mantissa[31]), .S(o_mantissa[47]), 
      .Z(n_30));
   MUX2_X1 i_1_102 (.A(o_mantissa[31]), .B(o_mantissa[32]), .S(o_mantissa[47]), 
      .Z(n_31));
   MUX2_X1 i_1_103 (.A(o_mantissa[32]), .B(o_mantissa[33]), .S(o_mantissa[47]), 
      .Z(n_32));
   MUX2_X1 i_1_104 (.A(o_mantissa[33]), .B(o_mantissa[34]), .S(o_mantissa[47]), 
      .Z(n_33));
   MUX2_X1 i_1_105 (.A(o_mantissa[34]), .B(o_mantissa[35]), .S(o_mantissa[47]), 
      .Z(n_34));
   MUX2_X1 i_1_106 (.A(o_mantissa[35]), .B(o_mantissa[36]), .S(o_mantissa[47]), 
      .Z(n_35));
   MUX2_X1 i_1_107 (.A(o_mantissa[36]), .B(o_mantissa[37]), .S(o_mantissa[47]), 
      .Z(n_36));
   MUX2_X1 i_1_108 (.A(o_mantissa[37]), .B(o_mantissa[38]), .S(o_mantissa[47]), 
      .Z(n_37));
   MUX2_X1 i_1_109 (.A(o_mantissa[38]), .B(o_mantissa[39]), .S(o_mantissa[47]), 
      .Z(n_38));
   MUX2_X1 i_1_110 (.A(o_mantissa[39]), .B(o_mantissa[40]), .S(o_mantissa[47]), 
      .Z(n_39));
   MUX2_X1 i_1_111 (.A(o_mantissa[40]), .B(o_mantissa[41]), .S(o_mantissa[47]), 
      .Z(n_40));
   MUX2_X1 i_1_112 (.A(o_mantissa[41]), .B(o_mantissa[42]), .S(o_mantissa[47]), 
      .Z(n_41));
   MUX2_X1 i_1_113 (.A(o_mantissa[42]), .B(o_mantissa[43]), .S(o_mantissa[47]), 
      .Z(n_42));
   MUX2_X1 i_1_114 (.A(o_mantissa[43]), .B(o_mantissa[44]), .S(o_mantissa[47]), 
      .Z(n_43));
   MUX2_X1 i_1_115 (.A(o_mantissa[44]), .B(o_mantissa[45]), .S(o_mantissa[47]), 
      .Z(n_44));
   MUX2_X1 i_1_116 (.A(o_mantissa[45]), .B(o_mantissa[46]), .S(o_mantissa[47]), 
      .Z(n_45));
   INV_X1 i_1_117 (.A(n_1_30), .ZN(n_1_74));
   INV_X1 i_1_118 (.A(n_1_29), .ZN(n_1_75));
   INV_X1 i_1_119 (.A(n_1_28), .ZN(n_1_76));
   INV_X1 i_1_120 (.A(n_1_27), .ZN(n_1_77));
   INV_X1 i_1_121 (.A(n_1_26), .ZN(n_1_78));
   INV_X1 i_1_122 (.A(n_1_25), .ZN(n_1_79));
   INV_X1 i_1_123 (.A(n_1_24), .ZN(n_1_80));
   INV_X1 i_1_84 (.A(n_1_15), .ZN(n_1_81));
   INV_X1 i_1_85 (.A(n_0), .ZN(n_1_82));
   INV_X1 i_1_126 (.A(n_1), .ZN(n_1_83));
   INV_X1 i_1_127 (.A(n_2), .ZN(n_1_84));
   INV_X1 i_1_128 (.A(n_3), .ZN(n_1_85));
   INV_X1 i_1_129 (.A(n_4), .ZN(n_1_86));
   INV_X1 i_1_130 (.A(n_5), .ZN(n_1_87));
   INV_X1 i_1_131 (.A(n_6), .ZN(n_1_88));
   INV_X1 i_1_132 (.A(n_7), .ZN(n_1_89));
   INV_X1 i_1_133 (.A(n_8), .ZN(n_1_90));
   INV_X1 i_1_134 (.A(n_9), .ZN(n_1_91));
   INV_X1 i_1_135 (.A(n_10), .ZN(n_1_92));
   INV_X1 i_1_136 (.A(n_11), .ZN(n_1_93));
   INV_X1 i_1_137 (.A(n_12), .ZN(n_1_94));
   INV_X1 i_1_138 (.A(n_13), .ZN(n_1_95));
   INV_X1 i_1_139 (.A(n_14), .ZN(n_1_96));
   INV_X1 i_1_140 (.A(n_15), .ZN(n_1_97));
   INV_X1 i_1_141 (.A(n_16), .ZN(n_1_98));
   INV_X1 i_1_142 (.A(n_17), .ZN(n_1_99));
   INV_X1 i_1_143 (.A(n_18), .ZN(n_1_100));
   INV_X1 i_1_144 (.A(n_19), .ZN(n_1_101));
   INV_X1 i_1_145 (.A(n_20), .ZN(n_1_102));
   INV_X1 i_1_146 (.A(n_21), .ZN(n_1_103));
   INV_X1 i_1_147 (.A(n_22), .ZN(n_1_104));
   INV_X1 i_1_86 (.A(n_1_65), .ZN(n_46));
   OAI222_X1 i_1_87 (.A1(n_1_105), .A2(o_mantissa[23]), .B1(o_mantissa[47]), 
      .B2(o_mantissa[22]), .C1(n_1_71), .C2(n_1_66), .ZN(n_1_65));
   NAND4_X1 i_1_88 (.A1(n_1_70), .A2(n_1_69), .A3(n_1_68), .A4(n_1_67), .ZN(
      n_1_66));
   NOR4_X1 i_1_89 (.A1(o_mantissa[6]), .A2(o_mantissa[5]), .A3(o_mantissa[4]), 
      .A4(o_mantissa[3]), .ZN(n_1_67));
   NOR3_X1 i_1_90 (.A1(o_mantissa[2]), .A2(o_mantissa[1]), .A3(o_mantissa[0]), 
      .ZN(n_1_68));
   NOR4_X1 i_1_91 (.A1(o_mantissa[14]), .A2(o_mantissa[13]), .A3(o_mantissa[12]), 
      .A4(o_mantissa[11]), .ZN(n_1_69));
   NOR4_X1 i_1_92 (.A1(o_mantissa[10]), .A2(o_mantissa[9]), .A3(o_mantissa[8]), 
      .A4(o_mantissa[7]), .ZN(n_1_70));
   NAND2_X1 i_1_93 (.A1(n_1_73), .A2(n_1_72), .ZN(n_1_71));
   NOR4_X1 i_1_124 (.A1(o_mantissa[22]), .A2(o_mantissa[19]), .A3(o_mantissa[17]), 
      .A4(o_mantissa[16]), .ZN(n_1_72));
   NOR4_X1 i_1_125 (.A1(o_mantissa[21]), .A2(o_mantissa[20]), .A3(o_mantissa[18]), 
      .A4(o_mantissa[15]), .ZN(n_1_73));
   INV_X1 i_1_148 (.A(o_mantissa[47]), .ZN(n_1_105));
endmodule

module registerNbits(clk, reset, en, inp, out);
   input clk;
   input reset;
   input en;
   input [31:0]inp;
   output [31:0]out;

   wire n_0_0;

   CLKGATETST_X1 clk_gate_out_reg (.CK(clk), .E(n_1), .SE(1'b0), .GCK(n_0));
   DFF_X1 \out_reg[31]  (.D(n_33), .CK(n_0), .Q(out[31]), .QN());
   DFF_X1 \out_reg[30]  (.D(n_32), .CK(n_0), .Q(out[30]), .QN());
   DFF_X1 \out_reg[29]  (.D(n_31), .CK(n_0), .Q(out[29]), .QN());
   DFF_X1 \out_reg[28]  (.D(n_30), .CK(n_0), .Q(out[28]), .QN());
   DFF_X1 \out_reg[27]  (.D(n_29), .CK(n_0), .Q(out[27]), .QN());
   DFF_X1 \out_reg[26]  (.D(n_28), .CK(n_0), .Q(out[26]), .QN());
   DFF_X1 \out_reg[25]  (.D(n_27), .CK(n_0), .Q(out[25]), .QN());
   DFF_X1 \out_reg[24]  (.D(n_26), .CK(n_0), .Q(out[24]), .QN());
   DFF_X1 \out_reg[23]  (.D(n_25), .CK(n_0), .Q(out[23]), .QN());
   DFF_X1 \out_reg[22]  (.D(n_24), .CK(n_0), .Q(out[22]), .QN());
   DFF_X1 \out_reg[21]  (.D(n_23), .CK(n_0), .Q(out[21]), .QN());
   DFF_X1 \out_reg[20]  (.D(n_22), .CK(n_0), .Q(out[20]), .QN());
   DFF_X1 \out_reg[19]  (.D(n_21), .CK(n_0), .Q(out[19]), .QN());
   DFF_X1 \out_reg[18]  (.D(n_20), .CK(n_0), .Q(out[18]), .QN());
   DFF_X1 \out_reg[17]  (.D(n_19), .CK(n_0), .Q(out[17]), .QN());
   DFF_X1 \out_reg[16]  (.D(n_18), .CK(n_0), .Q(out[16]), .QN());
   DFF_X1 \out_reg[15]  (.D(n_17), .CK(n_0), .Q(out[15]), .QN());
   DFF_X1 \out_reg[14]  (.D(n_16), .CK(n_0), .Q(out[14]), .QN());
   DFF_X1 \out_reg[13]  (.D(n_15), .CK(n_0), .Q(out[13]), .QN());
   DFF_X1 \out_reg[12]  (.D(n_14), .CK(n_0), .Q(out[12]), .QN());
   DFF_X1 \out_reg[11]  (.D(n_13), .CK(n_0), .Q(out[11]), .QN());
   DFF_X1 \out_reg[10]  (.D(n_12), .CK(n_0), .Q(out[10]), .QN());
   DFF_X1 \out_reg[9]  (.D(n_11), .CK(n_0), .Q(out[9]), .QN());
   DFF_X1 \out_reg[8]  (.D(n_10), .CK(n_0), .Q(out[8]), .QN());
   DFF_X1 \out_reg[7]  (.D(n_9), .CK(n_0), .Q(out[7]), .QN());
   DFF_X1 \out_reg[6]  (.D(n_8), .CK(n_0), .Q(out[6]), .QN());
   DFF_X1 \out_reg[5]  (.D(n_7), .CK(n_0), .Q(out[5]), .QN());
   DFF_X1 \out_reg[4]  (.D(n_6), .CK(n_0), .Q(out[4]), .QN());
   DFF_X1 \out_reg[3]  (.D(n_5), .CK(n_0), .Q(out[3]), .QN());
   DFF_X1 \out_reg[2]  (.D(n_4), .CK(n_0), .Q(out[2]), .QN());
   DFF_X1 \out_reg[1]  (.D(n_3), .CK(n_0), .Q(out[1]), .QN());
   DFF_X1 \out_reg[0]  (.D(n_2), .CK(n_0), .Q(out[0]), .QN());
   OR2_X1 i_0_0 (.A1(en), .A2(reset), .ZN(n_1));
   INV_X1 i_0_1 (.A(reset), .ZN(n_0_0));
   AND2_X1 i_0_2 (.A1(n_0_0), .A2(inp[0]), .ZN(n_2));
   AND2_X1 i_0_3 (.A1(n_0_0), .A2(inp[1]), .ZN(n_3));
   AND2_X1 i_0_4 (.A1(n_0_0), .A2(inp[2]), .ZN(n_4));
   AND2_X1 i_0_5 (.A1(n_0_0), .A2(inp[3]), .ZN(n_5));
   AND2_X1 i_0_6 (.A1(n_0_0), .A2(inp[4]), .ZN(n_6));
   AND2_X1 i_0_7 (.A1(n_0_0), .A2(inp[5]), .ZN(n_7));
   AND2_X1 i_0_8 (.A1(n_0_0), .A2(inp[6]), .ZN(n_8));
   AND2_X1 i_0_9 (.A1(n_0_0), .A2(inp[7]), .ZN(n_9));
   AND2_X1 i_0_10 (.A1(n_0_0), .A2(inp[8]), .ZN(n_10));
   AND2_X1 i_0_11 (.A1(n_0_0), .A2(inp[9]), .ZN(n_11));
   AND2_X1 i_0_12 (.A1(n_0_0), .A2(inp[10]), .ZN(n_12));
   AND2_X1 i_0_13 (.A1(n_0_0), .A2(inp[11]), .ZN(n_13));
   AND2_X1 i_0_14 (.A1(n_0_0), .A2(inp[12]), .ZN(n_14));
   AND2_X1 i_0_15 (.A1(n_0_0), .A2(inp[13]), .ZN(n_15));
   AND2_X1 i_0_16 (.A1(n_0_0), .A2(inp[14]), .ZN(n_16));
   AND2_X1 i_0_17 (.A1(n_0_0), .A2(inp[15]), .ZN(n_17));
   AND2_X1 i_0_18 (.A1(n_0_0), .A2(inp[16]), .ZN(n_18));
   AND2_X1 i_0_19 (.A1(n_0_0), .A2(inp[17]), .ZN(n_19));
   AND2_X1 i_0_20 (.A1(n_0_0), .A2(inp[18]), .ZN(n_20));
   AND2_X1 i_0_21 (.A1(n_0_0), .A2(inp[19]), .ZN(n_21));
   AND2_X1 i_0_22 (.A1(n_0_0), .A2(inp[20]), .ZN(n_22));
   AND2_X1 i_0_23 (.A1(n_0_0), .A2(inp[21]), .ZN(n_23));
   AND2_X1 i_0_24 (.A1(n_0_0), .A2(inp[22]), .ZN(n_24));
   AND2_X1 i_0_25 (.A1(n_0_0), .A2(inp[23]), .ZN(n_25));
   AND2_X1 i_0_26 (.A1(n_0_0), .A2(inp[24]), .ZN(n_26));
   AND2_X1 i_0_27 (.A1(n_0_0), .A2(inp[25]), .ZN(n_27));
   AND2_X1 i_0_28 (.A1(n_0_0), .A2(inp[26]), .ZN(n_28));
   AND2_X1 i_0_29 (.A1(n_0_0), .A2(inp[27]), .ZN(n_29));
   AND2_X1 i_0_30 (.A1(n_0_0), .A2(inp[28]), .ZN(n_30));
   AND2_X1 i_0_31 (.A1(n_0_0), .A2(inp[29]), .ZN(n_31));
   AND2_X1 i_0_32 (.A1(n_0_0), .A2(inp[30]), .ZN(n_32));
   AND2_X1 i_0_33 (.A1(n_0_0), .A2(inp[31]), .ZN(n_33));
endmodule

module FloatingPointMultiplierSingle(clk, reset, en, inputA, inputB, result, OF);
   input clk;
   input reset;
   input en;
   input [31:0]inputA;
   input [31:0]inputB;
   output [31:0]result;
   output OF;

   wire [31:0]A_reg;
   wire [31:0]B_reg;
   wire [31:0]out;

   registerNbits__0_18 regA (.clk(clk), .reset(reset), .en(en), .inp(inputA), 
      .out(A_reg));
   registerNbits__0_21 regB (.clk(clk), .reset(reset), .en(en), .inp(inputB), 
      .out(B_reg));
   FloatingPointMultiplier FloatingPointMultiplier_dut (.A(A_reg), .B(B_reg), 
      .O(out), .OF(OF));
   registerNbits outReg (.clk(clk), .reset(reset), .en(en), .inp(out), .out(
      result));
endmodule
