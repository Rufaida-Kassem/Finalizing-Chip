* SPICE NETLIST
***************************************

.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q 6
** N=21 EP=6 IP=0 FDC=28
M0 VSS 10 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 18 9 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 8 7 18 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 19 10 8 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 19 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 9 8 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 10 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 20 8 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 11 7 20 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 21 10 11 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 13 21 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 13 11 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 11 QN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 13 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 10 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 14 9 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 8 10 14 VDD PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 15 7 8 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 15 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 9 8 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 16 8 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 11 10 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 17 7 11 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 13 17 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 13 11 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 11 QN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_6
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6
** N=8 EP=6 IP=0 FDC=6
M0 8 A1 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5
** N=5 EP=5 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222_X1 C2 C1 VDD B1 B2 A2 VSS A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 13 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=675 $Y=90 $D=1
M3 VSS B2 13 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=865 $Y=90 $D=1
M4 14 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1055 $Y=90 $D=1
M5 ZN A1 14 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1245 $Y=90 $D=1
M6 10 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD C1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 10 B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=675 $Y=680 $D=0
M9 11 B2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=865 $Y=680 $D=0
M10 ZN A2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1055 $Y=680 $D=0
M11 11 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1245 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DLH_X1 G Q D VSS VDD
** N=13 EP=5 IP=0 FDC=16
M0 VSS G 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07 $X=170 $Y=90 $D=1
M1 Q 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS 6 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=755 $Y=215 $D=1
M3 12 D VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=945 $Y=215 $D=1
M4 8 7 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1135 $Y=215 $D=1
M5 13 6 8 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=1325 $Y=335 $D=1
M6 VSS 9 13 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=335 $D=1
M7 9 8 VSS VSS NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=335 $D=1
M8 VDD G 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=170 $Y=995 $D=0
M9 Q 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M10 VDD 6 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=755 $Y=815 $D=0
M11 10 D VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=945 $Y=815 $D=0
M12 8 6 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1135 $Y=815 $D=0
M13 11 7 8 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=1325 $Y=1040 $D=0
M14 VDD 9 11 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=1040 $D=0
M15 9 8 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=1040 $D=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 8 A3 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 9 A1 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 11 A3 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 9 A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR4_X2 A1 A2 A3 ZN A4 VSS VDD
** N=13 EP=7 IP=0 FDC=16
M0 ZN A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A3 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=945 $Y=90 $D=1
M5 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1135 $Y=90 $D=1
M6 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1325 $Y=90 $D=1
M7 VSS A4 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1515 $Y=90 $D=1
M8 8 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 9 A3 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 10 A2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 ZN A1 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
M12 11 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=945 $Y=680 $D=0
M13 12 A2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1135 $Y=680 $D=0
M14 13 A3 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1325 $Y=680 $D=0
M15 VDD A4 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1515 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 8 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 7 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 VSS B2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS
** N=10 EP=7 IP=0 FDC=8
M0 9 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 8 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 8 A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 5 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD
** N=10 EP=7 IP=0 FDC=8
M0 VSS B2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 8 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 8 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 10 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 11 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7
** N=9 EP=7 IP=0 FDC=6
M0 ZN B2 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 8 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 8 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD
** N=6 EP=5 IP=0 FDC=4
M0 6 A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS
** N=6 EP=5 IP=0 FDC=4
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT INV_X2 A ZN VSS VDD
** N=4 EP=4 IP=0 FDC=4
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143
** N=261 EP=143 IP=4135 FDC=2080
X2159 243 18 68 67 158 68 DFF_X1 $T=18100 68200 1 0 $X=17985 $Y=66685
X2160 244 18 68 67 160 68 DFF_X1 $T=21330 68200 1 0 $X=21215 $Y=66685
X2161 159 26 68 67 161 68 DFF_X1 $T=22280 65400 0 0 $X=22165 $Y=65285
X2162 237 26 68 67 163 68 DFF_X1 $T=28740 65400 1 180 $X=25395 $Y=65285
X2163 224 18 68 67 162 68 DFF_X1 $T=26080 68200 0 0 $X=25965 $Y=68085
X2164 225 26 68 67 164 68 DFF_X1 $T=28550 65400 1 0 $X=28435 $Y=63885
X2165 245 18 68 67 29 68 DFF_X1 $T=30640 68200 0 0 $X=30525 $Y=68085
X2166 246 18 68 67 40 68 DFF_X1 $T=34630 65400 0 0 $X=34515 $Y=65285
X2167 227 26 68 67 87 68 DFF_X1 $T=37860 65400 0 0 $X=37745 $Y=65285
X2168 247 18 68 67 53 68 DFF_X1 $T=38620 68200 1 0 $X=38505 $Y=66685
X2169 248 26 68 67 113 68 DFF_X1 $T=41660 65400 1 0 $X=41545 $Y=63885
X2170 249 18 68 67 47 68 DFF_X1 $T=42230 68200 1 0 $X=42115 $Y=66685
X2171 259 18 68 67 42 68 DFF_X1 $T=45460 68200 1 180 $X=42115 $Y=68085
X2172 167 26 68 67 88 68 DFF_X1 $T=44320 62600 0 0 $X=44205 $Y=62485
X2173 260 26 68 67 103 68 DFF_X1 $T=48120 65400 0 180 $X=44775 $Y=63885
X2174 250 18 68 67 39 68 DFF_X1 $T=45460 68200 1 0 $X=45345 $Y=66685
X2175 168 18 68 67 114 68 DFF_X1 $T=46790 62600 1 0 $X=46675 $Y=61085
X2176 229 18 68 67 46 68 DFF_X1 $T=52300 62600 0 0 $X=52185 $Y=62485
X2177 238 18 68 67 37 68 DFF_X1 $T=57810 62600 0 180 $X=54465 $Y=61085
X2178 230 18 68 67 165 68 DFF_X1 $T=54770 65400 0 0 $X=54655 $Y=65285
X2179 239 26 68 67 61 68 DFF_X1 $T=55530 62600 0 0 $X=55415 $Y=62485
X2180 251 18 68 67 166 68 DFF_X1 $T=55530 68200 0 0 $X=55415 $Y=68085
X2181 195 26 68 67 60 68 DFF_X1 $T=58760 62600 0 0 $X=58645 $Y=62485
X2182 252 26 68 67 49 68 DFF_X1 $T=58760 65400 1 0 $X=58645 $Y=63885
X2183 242 65 68 67 128 68 DFF_X1 $T=58760 68200 1 0 $X=58645 $Y=66685
X2184 194 65 68 67 129 68 DFF_X1 $T=58760 68200 0 0 $X=58645 $Y=68085
X2185 197 65 68 67 92 68 DFF_X1 $T=59710 62600 1 0 $X=59595 $Y=61085
X2186 131 65 68 67 130 68 DFF_X1 $T=62370 59800 0 0 $X=62255 $Y=59685
X2187 214 65 68 67 91 68 DFF_X1 $T=62370 68200 0 0 $X=62255 $Y=68085
X2188 232 65 68 67 105 68 DFF_X1 $T=65790 62600 1 0 $X=65675 $Y=61085
X2189 215 65 68 67 106 68 DFF_X1 $T=65790 65400 0 0 $X=65675 $Y=65285
X2190 196 65 68 67 124 68 DFF_X1 $T=66170 59800 0 0 $X=66055 $Y=59685
X2191 253 65 68 67 116 68 DFF_X1 $T=66170 65400 1 0 $X=66055 $Y=63885
X2287 86 15 68 67 256 68 AND2_X1 $T=17530 68200 0 0 $X=17415 $Y=68085
X2288 86 21 68 67 213 68 AND2_X1 $T=21140 68200 0 0 $X=21025 $Y=68085
X2289 84 24 68 67 159 68 AND2_X1 $T=23990 68200 1 180 $X=23115 $Y=68085
X2290 86 28 68 67 224 68 AND2_X1 $T=25320 68200 0 0 $X=25205 $Y=68085
X2291 84 30 68 67 237 68 AND2_X1 $T=27790 68200 0 180 $X=26915 $Y=66685
X2292 84 31 68 67 225 68 AND2_X1 $T=29310 68200 0 0 $X=29195 $Y=68085
X2293 86 32 68 67 245 68 AND2_X1 $T=30640 68200 1 0 $X=30525 $Y=66685
X2294 86 36 68 67 246 68 AND2_X1 $T=34630 68200 1 180 $X=33755 $Y=68085
X2295 86 38 68 67 247 68 AND2_X1 $T=36340 68200 0 0 $X=36225 $Y=68085
X2296 84 41 68 67 227 68 AND2_X1 $T=39570 68200 1 180 $X=38695 $Y=68085
X2297 86 43 68 67 112 68 AND2_X1 $T=40900 65400 1 0 $X=40785 $Y=63885
X2298 84 44 68 67 248 68 AND2_X1 $T=41090 65400 0 0 $X=40975 $Y=65285
X2299 86 45 68 67 249 68 AND2_X1 $T=41090 68200 0 0 $X=40975 $Y=68085
X2300 84 48 68 67 167 68 AND2_X1 $T=45270 65400 1 180 $X=44395 $Y=65285
X2301 86 50 68 67 259 68 AND2_X1 $T=46220 68200 1 180 $X=45345 $Y=68085
X2302 84 51 68 67 260 68 AND2_X1 $T=47170 65400 1 180 $X=46295 $Y=65285
X2303 90 169 68 67 242 68 AND2_X1 $T=49260 65400 0 0 $X=49145 $Y=65285
X2304 86 52 68 67 250 68 AND2_X1 $T=50020 68200 1 180 $X=49145 $Y=68085
X2305 86 54 68 67 168 68 AND2_X1 $T=50780 65400 1 180 $X=49905 $Y=65285
X2306 86 55 68 67 229 68 AND2_X1 $T=50780 65400 0 0 $X=50665 $Y=65285
X2307 86 56 68 67 230 68 AND2_X1 $T=52490 68200 1 180 $X=51615 $Y=68085
X2308 86 57 68 67 238 68 AND2_X1 $T=52110 65400 1 0 $X=51995 $Y=63885
X2309 86 58 68 67 251 68 AND2_X1 $T=52490 68200 0 0 $X=52375 $Y=68085
X2310 84 59 68 67 239 68 AND2_X1 $T=54200 65400 1 0 $X=54085 $Y=63885
X2311 90 170 68 67 194 68 AND2_X1 $T=56290 65400 1 0 $X=56175 $Y=63885
X2312 84 62 68 67 252 68 AND2_X1 $T=58000 65400 0 0 $X=57885 $Y=65285
X2313 84 64 68 67 195 68 AND2_X1 $T=58760 65400 0 0 $X=58645 $Y=65285
X2314 90 171 68 67 196 68 AND2_X1 $T=59520 59800 0 0 $X=59405 $Y=59685
X2315 90 172 68 67 214 68 AND2_X1 $T=62370 65400 0 0 $X=62255 $Y=65285
X2316 90 173 68 67 232 68 AND2_X1 $T=63130 62600 1 0 $X=63015 $Y=61085
X2317 90 174 68 67 215 68 AND2_X1 $T=63130 65400 0 0 $X=63015 $Y=65285
X2318 90 175 68 67 253 68 AND2_X1 $T=63510 62600 0 0 $X=63395 $Y=62485
X2319 90 176 68 67 197 68 AND2_X1 $T=63890 65400 0 0 $X=63775 $Y=65285
X2536 137 68 67 68 68 INV_X1 $T=1760 59800 0 0 $X=1645 $Y=59685
X2537 240 68 67 199 68 INV_X1 $T=5180 62600 1 180 $X=4685 $Y=62485
X2538 3 68 67 2 68 INV_X1 $T=6320 65400 0 180 $X=5825 $Y=63885
X2539 138 68 67 180 68 INV_X1 $T=8220 59800 1 180 $X=7725 $Y=59685
X2540 201 68 67 254 68 INV_X1 $T=8600 65400 1 180 $X=8105 $Y=65285
X2541 218 68 67 183 68 INV_X1 $T=8600 65400 0 0 $X=8485 $Y=65285
X2542 146 68 67 241 68 INV_X1 $T=12400 65400 0 180 $X=11905 $Y=63885
X2543 185 68 67 221 68 INV_X1 $T=14110 65400 0 0 $X=13995 $Y=65285
X2544 79 68 67 149 68 INV_X1 $T=14870 62600 0 0 $X=14755 $Y=62485
X2545 222 68 67 209 68 INV_X1 $T=16200 65400 0 180 $X=15705 $Y=63885
X2546 226 68 67 169 68 INV_X1 $T=38430 65400 1 0 $X=38315 $Y=63885
X2547 193 68 67 174 68 INV_X1 $T=43940 62600 0 0 $X=43825 $Y=62485
X2548 228 68 67 175 68 INV_X1 $T=46410 62600 1 0 $X=46295 $Y=61085
X2549 115 68 67 170 68 INV_X1 $T=55910 65400 1 0 $X=55795 $Y=63885
X2550 63 68 67 171 68 INV_X1 $T=58760 59800 0 0 $X=58645 $Y=59685
X2551 141 68 67 173 68 INV_X1 $T=59140 59800 0 0 $X=59025 $Y=59685
X2552 231 68 67 172 68 INV_X1 $T=59710 62600 0 180 $X=59215 $Y=61085
X2553 261 68 67 176 68 INV_X1 $T=62370 62600 0 0 $X=62255 $Y=62485
X2629 14 9 67 8 7 125 68 77 186 AOI222_X1 $T=15060 62600 0 180 $X=13425 $Y=61085
X2630 125 10 67 11 14 7 68 80 205 AOI222_X1 $T=15060 62600 1 0 $X=14945 $Y=61085
X2631 125 12 67 13 7 14 68 97 222 AOI222_X1 $T=15440 59800 0 0 $X=15325 $Y=59685
X2632 35 161 67 34 158 33 68 139 226 AOI222_X1 $T=32160 62600 1 180 $X=30525 $Y=62485
X2633 35 163 67 34 160 33 68 120 193 AOI222_X1 $T=33870 62600 0 180 $X=32235 $Y=61085
X2634 35 164 67 34 162 33 68 121 228 AOI222_X1 $T=33870 62600 1 0 $X=33755 $Y=61085
X2635 35 113 67 34 53 33 68 127 89 AOI222_X1 $T=50780 59800 1 180 $X=49145 $Y=59685
X2636 35 60 67 34 165 33 68 140 261 AOI222_X1 $T=57240 59800 0 0 $X=57125 $Y=59685
X2637 35 61 67 34 166 33 68 123 231 AOI222_X1 $T=57810 62600 1 0 $X=57695 $Y=61085
X2647 101 80 158 68 67 DLH_X1 $T=24180 62600 1 180 $X=22165 $Y=62485
X2648 101 13 160 68 67 DLH_X1 $T=24180 62600 0 0 $X=24065 $Y=62485
X2649 101 136 161 68 67 DLH_X1 $T=25320 62600 1 0 $X=25205 $Y=61085
X2650 101 118 29 68 67 DLH_X1 $T=25700 59800 0 0 $X=25585 $Y=59685
X2651 101 8 162 68 67 DLH_X1 $T=26650 65400 1 0 $X=26535 $Y=63885
X2652 101 85 163 68 67 DLH_X1 $T=27220 62600 1 0 $X=27105 $Y=61085
X2653 101 119 164 68 67 DLH_X1 $T=29500 59800 0 0 $X=29385 $Y=59685
X2654 33 110 37 68 67 DLH_X1 $T=34060 59800 0 0 $X=33945 $Y=59685
X2655 33 27 165 68 67 DLH_X1 $T=35960 59800 0 0 $X=35845 $Y=59685
X2656 33 11 39 68 67 DLH_X1 $T=35960 62600 0 0 $X=35845 $Y=62485
X2657 33 9 40 68 67 DLH_X1 $T=36530 65400 1 0 $X=36415 $Y=63885
X2658 33 23 166 68 67 DLH_X1 $T=39950 62600 0 180 $X=37935 $Y=61085
X2659 33 10 42 68 67 DLH_X1 $T=39950 62600 1 0 $X=39835 $Y=61085
X2660 33 12 53 68 67 DLH_X1 $T=39950 62600 0 0 $X=39835 $Y=62485
X2661 33 102 46 68 67 DLH_X1 $T=41090 59800 0 0 $X=40975 $Y=59685
X2662 33 77 47 68 67 DLH_X1 $T=44130 62600 0 180 $X=42115 $Y=61085
X2663 33 122 103 68 67 DLH_X1 $T=42990 59800 0 0 $X=42875 $Y=59685
X2664 33 104 49 68 67 DLH_X1 $T=44890 59800 0 0 $X=44775 $Y=59685
X2665 166 165 39 40 68 67 111 OR4_X1 $T=39000 59800 1 180 $X=37745 $Y=59685
X2666 87 67 164 163 161 67 68 NOR4_X1 $T=31400 62600 0 180 $X=30335 $Y=61085
X2667 158 160 162 109 29 68 67 NOR4_X2 $T=28930 62600 0 0 $X=28815 $Y=62485
X2680 68 1 216 233 68 67 AOI21_X1 $T=2330 68200 1 0 $X=2215 $Y=66685
X2681 254 1 210 203 68 67 AOI21_X1 $T=9360 68200 0 0 $X=9245 $Y=68085
X2682 241 1 235 76 68 67 AOI21_X1 $T=11830 65400 0 0 $X=11715 $Y=65285
X2683 221 1 187 208 68 67 AOI21_X1 $T=14490 65400 0 0 $X=14375 $Y=65285
X2684 190 19 99 211 68 67 AOI21_X1 $T=19430 62600 1 0 $X=19315 $Y=61085
X2685 25 23 126 258 68 67 AOI21_X1 $T=23800 62600 0 180 $X=22925 $Y=61085
X2686 25 11 143 257 68 67 AOI21_X1 $T=23800 62600 1 0 $X=23685 $Y=61085
X2687 25 9 100 223 68 67 AOI21_X1 $T=25320 62600 0 180 $X=24445 $Y=61085
X2688 25 27 117 236 68 67 AOI21_X1 $T=24940 59800 0 0 $X=24825 $Y=59685
X2691 186 3 68 5 4 67 2 207 OAI221_X1 $T=13540 62600 1 180 $X=12285 $Y=62485
X2692 75 6 68 147 148 67 16 78 OAI221_X1 $T=13350 59800 0 0 $X=13235 $Y=59685
X2693 81 6 68 151 152 67 16 107 OAI221_X1 $T=17340 65400 0 0 $X=17225 $Y=65285
X2694 98 6 68 153 154 67 16 134 OAI221_X1 $T=17910 59800 0 0 $X=17795 $Y=59685
X2695 189 16 68 150 17 67 6 258 OAI221_X1 $T=18290 62600 0 0 $X=18175 $Y=62485
X2696 191 16 68 155 20 67 6 236 OAI221_X1 $T=19620 65400 1 0 $X=19505 $Y=63885
X2697 108 6 68 156 157 67 16 257 OAI221_X1 $T=20760 65400 1 0 $X=20645 $Y=63885
X2698 212 16 68 192 22 67 6 223 OAI221_X1 $T=21140 62600 1 0 $X=21025 $Y=61085
X2699 216 94 67 95 132 177 68 AOI22_X1 $T=2900 65400 0 180 $X=1835 $Y=63885
X2700 177 94 67 95 142 93 68 AOI22_X1 $T=3090 59800 1 180 $X=2025 $Y=59685
X2701 199 5 67 1 177 66 68 AOI22_X1 $T=3280 62600 1 180 $X=2215 $Y=62485
X2702 234 94 67 95 148 216 68 AOI22_X1 $T=4040 68200 0 180 $X=2975 $Y=66685
X2703 69 3 67 2 178 219 68 AOI22_X1 $T=4990 65400 1 0 $X=4875 $Y=63885
X2704 199 1 67 5 234 179 68 AOI22_X1 $T=4990 65400 0 0 $X=4875 $Y=65285
X2705 234 95 67 94 152 145 68 AOI22_X1 $T=4990 68200 0 0 $X=4875 $Y=68085
X2706 70 8 67 2 66 180 68 AOI22_X1 $T=5180 59800 0 0 $X=5065 $Y=59685
X2707 71 3 67 2 240 181 68 AOI22_X1 $T=5370 62600 1 0 $X=5255 $Y=61085
X2708 254 5 67 1 200 179 68 AOI22_X1 $T=6890 65400 0 0 $X=6775 $Y=65285
X2709 200 94 67 95 189 145 68 AOI22_X1 $T=7460 68200 1 0 $X=7345 $Y=66685
X2710 181 3 67 2 201 74 68 AOI22_X1 $T=7650 62600 0 0 $X=7535 $Y=62485
X2711 125 80 67 10 181 14 68 AOI22_X1 $T=9360 62600 0 180 $X=8295 $Y=61085
X2712 125 13 67 12 219 14 68 AOI22_X1 $T=9360 62600 1 0 $X=9245 $Y=61085
X2713 183 1 67 5 204 184 68 AOI22_X1 $T=9930 65400 0 0 $X=9815 $Y=65285
X2714 125 8 67 77 182 14 68 AOI22_X1 $T=10310 62600 1 0 $X=10195 $Y=61085
X2715 210 94 67 95 73 204 68 AOI22_X1 $T=10690 68200 0 0 $X=10575 $Y=68085
X2716 204 94 67 95 154 200 68 AOI22_X1 $T=10880 65400 0 0 $X=10765 $Y=65285
X2717 182 3 67 2 255 4 68 AOI22_X1 $T=11070 65400 1 0 $X=10955 $Y=63885
X2718 75 82 67 19 147 148 68 AOI22_X1 $T=12210 59800 1 180 $X=11145 $Y=59685
X2719 74 3 67 2 146 205 68 AOI22_X1 $T=11450 62600 0 0 $X=11335 $Y=62485
X2720 184 1 67 5 220 221 68 AOI22_X1 $T=12400 68200 1 0 $X=12285 $Y=66685
X2721 235 207 67 95 212 187 68 AOI22_X1 $T=13730 65400 1 0 $X=13615 $Y=63885
X2722 133 2 67 3 185 72 68 AOI22_X1 $T=14490 59800 0 0 $X=14375 $Y=59685
X2723 220 95 67 94 157 188 68 AOI22_X1 $T=14490 68200 0 0 $X=14375 $Y=68085
X2724 187 94 67 95 190 188 68 AOI22_X1 $T=14680 68200 1 0 $X=14565 $Y=66685
X2725 220 94 67 95 191 210 68 AOI22_X1 $T=15440 68200 0 0 $X=15325 $Y=68085
X2726 81 82 67 19 151 152 68 AOI22_X1 $T=16390 65400 0 0 $X=16275 $Y=65285
X2727 154 19 67 82 153 98 68 AOI22_X1 $T=16960 59800 0 0 $X=16845 $Y=59685
X2728 189 19 67 82 150 17 68 AOI22_X1 $T=17340 62600 0 0 $X=17225 $Y=62485
X2729 20 82 67 19 155 191 68 AOI22_X1 $T=18480 65400 0 0 $X=18365 $Y=65285
X2730 83 82 67 97 135 25 68 AOI22_X1 $T=20950 59800 0 0 $X=20835 $Y=59685
X2731 22 82 67 19 192 212 68 AOI22_X1 $T=21900 62600 1 180 $X=20835 $Y=62485
X2732 108 82 67 19 156 157 68 AOI22_X1 $T=20950 65400 0 0 $X=20835 $Y=65285
X2733 256 68 67 243 CLKBUF_X1 $T=18290 68200 0 0 $X=18175 $Y=68085
X2734 213 68 67 244 CLKBUF_X1 $T=20570 68200 0 0 $X=20455 $Y=68085
X2735 72 3 68 218 2 96 67 OAI22_X1 $T=8790 59800 0 0 $X=8675 $Y=59685
X2736 83 6 68 211 16 190 67 OAI22_X1 $T=20380 62600 1 180 $X=19315 $Y=62485
X2739 209 2 67 1 149 68 3 208 AOI221_X1 $T=15820 65400 0 180 $X=14565 $Y=63885
X2740 183 1 145 198 68 67 68 OAI21_X1 $T=7460 68200 1 180 $X=6585 $Y=68085
X2741 180 2 179 217 68 67 68 OAI21_X1 $T=7460 65400 1 0 $X=7345 $Y=63885
X2742 149 3 184 202 68 67 68 OAI21_X1 $T=11070 65400 0 180 $X=10195 $Y=63885
X2743 241 1 188 206 68 67 68 OAI21_X1 $T=12970 68200 1 180 $X=12095 $Y=68085
X2744 178 68 1 198 67 NAND2_X1 $T=4420 68200 0 0 $X=4305 $Y=68085
X2745 182 68 2 217 67 NAND2_X1 $T=8790 65400 0 180 $X=8105 $Y=63885
X2746 219 68 3 202 67 NAND2_X1 $T=9740 65400 1 0 $X=9625 $Y=63885
X2747 255 68 1 206 67 NAND2_X1 $T=11640 68200 0 0 $X=11525 $Y=68085
X2748 178 67 1 233 68 NOR2_X1 $T=3470 68200 1 180 $X=2785 $Y=68085
X2749 255 67 1 203 68 NOR2_X1 $T=10690 68200 1 180 $X=10005 $Y=68085
X2750 5 1 68 67 INV_X2 $T=2330 68200 0 0 $X=2215 $Y=68085
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN
** N=8 EP=6 IP=0 FDC=6
M0 ZN A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 8 A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S
** N=19 EP=7 IP=0 FDC=28
M0 VSS 8 CO VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 17 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 8 A 17 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 9 CI 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 9 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 11 B VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 11 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 13 8 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 18 CI 13 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 19 B 18 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 19 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 13 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 8 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 14 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 8 A 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 10 CI 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 10 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 12 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 12 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 13 8 12 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 15 CI 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 16 B 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD
** N=9 EP=5 IP=0 FDC=10
M0 9 A 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 7 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 7 B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 6 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 8 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS
** N=10 EP=7 IP=0 FDC=8
M0 ZN C2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 8 C1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 10 A 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 9 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN
** N=14 EP=9 IP=0 FDC=12
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 10 B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 11 B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 11 A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 12 C2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 13 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 14 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI211_X1 C2 C1 B VSS A ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 10 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN C1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN C2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 8 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 9 B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD
** N=7 EP=5 IP=0 FDC=8
M0 ZN A2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 6 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 6 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 7 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 106 107 108 109 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
** N=358 EP=199 IP=4828 FDC=1748
M0 81 82 34 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=7075 $Y=53695 $D=1
M1 34 84 81 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7265 $Y=53695 $D=1
M2 81 4 34 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7455 $Y=53695 $D=1
M3 34 4 81 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7645 $Y=53695 $D=1
M4 81 84 34 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7835 $Y=53695 $D=1
M5 34 82 81 34 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=8025 $Y=53695 $D=1
M6 355 82 79 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=7075 $Y=52890 $D=0
M7 356 84 355 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7265 $Y=52890 $D=0
M8 81 4 356 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7455 $Y=52890 $D=0
M9 357 4 81 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7645 $Y=52890 $D=0
M10 358 84 357 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7835 $Y=52890 $D=0
M11 79 82 358 79 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=8025 $Y=52890 $D=0
X2326 171 69 34 79 140 34 DFF_X1 $T=54580 51400 0 0 $X=54465 $Y=51285
X2327 339 73 34 79 253 34 DFF_X1 $T=58760 57000 1 0 $X=58645 $Y=55485
X2328 323 73 34 79 254 34 DFF_X1 $T=59140 54200 1 0 $X=59025 $Y=52685
X2329 346 73 34 79 252 34 DFF_X1 $T=60470 57000 0 0 $X=60355 $Y=56885
X2330 338 77 34 79 185 34 DFF_X1 $T=65790 51400 0 0 $X=65675 $Y=51285
X2331 352 77 34 79 163 34 DFF_X1 $T=65790 57000 1 0 $X=65675 $Y=55485
X2332 297 77 34 79 143 34 DFF_X1 $T=65790 57000 0 0 $X=65675 $Y=56885
X2333 322 77 34 79 164 34 DFF_X1 $T=66170 54200 0 0 $X=66055 $Y=54085
X2383 4 5 34 79 15 34 AND2_X1 $T=9360 54200 1 180 $X=8485 $Y=54085
X2384 119 255 34 79 155 34 AND2_X1 $T=58950 51400 0 0 $X=58835 $Y=51285
X2385 119 256 34 79 297 34 AND2_X1 $T=59900 59800 0 180 $X=59025 $Y=58285
X2386 119 257 34 79 352 34 AND2_X1 $T=59710 57000 0 0 $X=59595 $Y=56885
X2387 119 258 34 79 184 34 AND2_X1 $T=61230 59800 1 0 $X=61115 $Y=58285
X2388 119 259 34 79 338 34 AND2_X1 $T=63130 51400 1 180 $X=62255 $Y=51285
X2389 119 260 34 79 322 34 AND2_X1 $T=63320 54200 1 0 $X=63205 $Y=52685
X2390 120 74 34 79 346 34 AND2_X1 $T=64460 59800 0 180 $X=63585 $Y=58285
X2391 120 75 34 79 323 34 AND2_X1 $T=64080 54200 1 0 $X=63965 $Y=52685
X2392 120 76 34 79 339 34 AND2_X1 $T=64080 57000 1 0 $X=63965 $Y=55485
X2917 347 34 79 121 34 INV_X1 $T=2710 54200 0 180 $X=2215 $Y=52685
X2918 26 34 79 27 34 INV_X1 $T=16200 54200 0 180 $X=15705 $Y=52685
X2919 218 34 79 268 34 INV_X1 $T=16200 54200 1 180 $X=15705 $Y=54085
X2920 307 34 79 304 34 INV_X1 $T=19430 54200 0 180 $X=18935 $Y=52685
X2921 354 34 79 305 34 INV_X1 $T=20760 54200 1 180 $X=20265 $Y=54085
X2922 353 34 79 273 34 INV_X1 $T=21140 54200 1 180 $X=20645 $Y=54085
X2923 310 34 79 276 34 INV_X1 $T=23230 51400 1 180 $X=22735 $Y=51285
X2924 342 34 79 327 34 INV_X1 $T=23610 57000 0 180 $X=23115 $Y=55485
X2925 277 34 79 221 34 INV_X1 $T=23990 57000 0 180 $X=23495 $Y=55485
X2926 343 34 79 308 34 INV_X1 $T=24180 57000 1 180 $X=23685 $Y=56885
X2927 30 34 79 227 34 INV_X1 $T=31400 54200 1 0 $X=31285 $Y=52685
X2928 42 34 79 283 34 INV_X1 $T=31400 54200 0 0 $X=31285 $Y=54085
X2929 21 34 79 228 34 INV_X1 $T=31590 57000 1 0 $X=31475 $Y=55485
X2930 39 34 79 314 34 INV_X1 $T=33110 54200 0 180 $X=32615 $Y=52685
X2931 11 34 79 234 34 INV_X1 $T=32730 57000 0 0 $X=32615 $Y=56885
X2932 223 34 79 282 34 INV_X1 $T=34440 54200 0 0 $X=34325 $Y=54085
X2933 44 34 79 231 34 INV_X1 $T=35200 57000 0 180 $X=34705 $Y=55485
X2934 19 34 79 233 34 INV_X1 $T=35200 59800 1 0 $X=35085 $Y=58285
X2935 10 34 79 235 34 INV_X1 $T=36910 59800 0 180 $X=36415 $Y=58285
X2936 8 34 79 284 34 INV_X1 $T=38240 54200 0 180 $X=37745 $Y=52685
X2937 225 34 79 241 34 INV_X1 $T=38050 54200 0 0 $X=37935 $Y=54085
X2938 50 34 79 238 34 INV_X1 $T=38240 57000 0 0 $X=38125 $Y=56885
X2939 41 34 79 239 34 INV_X1 $T=39570 54200 0 0 $X=39455 $Y=54085
X2940 51 34 79 285 34 INV_X1 $T=40140 57000 1 180 $X=39645 $Y=56885
X2941 32 34 79 286 34 INV_X1 $T=40900 57000 0 0 $X=40785 $Y=56885
X2942 36 34 79 244 34 INV_X1 $T=41850 54200 1 180 $X=41355 $Y=54085
X2943 320 34 79 255 34 INV_X1 $T=50590 54200 0 0 $X=50475 $Y=54085
X2944 189 34 79 295 34 INV_X1 $T=51730 54200 0 0 $X=51615 $Y=54085
X2945 118 34 79 296 34 INV_X1 $T=53820 54200 1 0 $X=53705 $Y=52685
X2946 193 34 79 335 34 INV_X1 $T=55150 54200 1 0 $X=55035 $Y=52685
X2947 70 34 79 139 34 INV_X1 $T=57050 54200 0 0 $X=56935 $Y=54085
X2948 190 34 79 170 34 INV_X1 $T=57430 54200 0 0 $X=57315 $Y=54085
X2949 141 34 79 336 34 INV_X1 $T=57810 51400 0 0 $X=57695 $Y=51285
X2950 191 34 79 337 34 INV_X1 $T=57810 54200 0 0 $X=57695 $Y=54085
X2951 192 34 79 256 34 INV_X1 $T=58000 59800 1 0 $X=57885 $Y=58285
X2952 294 34 79 257 34 INV_X1 $T=58380 57000 1 0 $X=58265 $Y=55485
X2953 351 34 79 260 34 INV_X1 $T=59330 54200 0 0 $X=59215 $Y=54085
X2954 321 34 79 258 34 INV_X1 $T=59330 57000 0 0 $X=59215 $Y=56885
X2955 142 34 79 259 34 INV_X1 $T=59710 51400 0 0 $X=59595 $Y=51285
X3070 17 10 79 12 14 15 34 78 194 AOI222_X1 $T=12590 57000 1 0 $X=12475 $Y=55485
X3071 17 11 79 13 14 15 34 16 198 AOI222_X1 $T=12590 57000 0 0 $X=12475 $Y=56885
X3072 17 19 79 20 14 15 34 92 166 AOI222_X1 $T=14110 57000 1 0 $X=13995 $Y=55485
X3073 14 18 79 21 17 15 34 91 90 AOI222_X1 $T=14110 57000 0 0 $X=13995 $Y=56885
X3074 14 25 79 32 17 15 34 88 89 AOI222_X1 $T=16960 59800 0 180 $X=15325 $Y=58285
X3075 99 223 79 35 37 38 34 49 224 AOI222_X1 $T=26840 54200 0 0 $X=26725 $Y=54085
X3076 38 225 79 40 37 99 34 104 348 AOI222_X1 $T=28360 54200 0 0 $X=28245 $Y=54085
X3077 38 41 79 226 99 37 34 103 220 AOI222_X1 $T=28740 54200 1 0 $X=28625 $Y=52685
X3078 332 242 79 244 41 51 34 286 237 AOI222_X1 $T=38810 57000 1 0 $X=38695 $Y=55485
X3079 111 43 79 52 53 54 34 112 320 AOI222_X1 $T=40330 59800 1 0 $X=40215 $Y=58285
X3080 111 61 79 52 63 54 34 116 294 AOI222_X1 $T=48310 57000 0 0 $X=48195 $Y=56885
X3081 111 67 79 52 60 54 34 295 65 AOI222_X1 $T=52680 59800 0 180 $X=51045 $Y=58285
X3082 111 62 79 52 68 54 34 296 169 AOI222_X1 $T=52680 59800 1 0 $X=52565 $Y=58285
X3083 111 253 79 52 165 54 34 335 321 AOI222_X1 $T=56860 57000 1 0 $X=56745 $Y=55485
X3084 111 254 79 52 140 54 34 336 351 AOI222_X1 $T=57620 54200 1 0 $X=57505 $Y=52685
X3085 111 252 79 52 72 54 34 337 162 AOI222_X1 $T=57810 57000 0 0 $X=57695 $Y=56885
X3101 182 183 43 34 79 DLH_X1 $T=30830 57000 0 0 $X=30715 $Y=56885
X3102 54 30 45 34 79 DLH_X1 $T=35200 59800 0 180 $X=33185 $Y=58285
X3103 54 226 57 34 79 DLH_X1 $T=42230 51400 0 0 $X=42115 $Y=51285
X3104 54 225 56 34 79 DLH_X1 $T=42230 57000 0 0 $X=42115 $Y=56885
X3105 54 49 61 34 79 DLH_X1 $T=44890 59800 1 0 $X=44775 $Y=58285
X3106 54 55 64 34 79 DLH_X1 $T=52490 57000 0 180 $X=50475 $Y=55485
X3107 54 44 252 34 79 DLH_X1 $T=52490 57000 1 0 $X=52375 $Y=55485
X3108 54 223 253 34 79 DLH_X1 $T=55150 54200 1 180 $X=53135 $Y=54085
X3109 54 48 254 34 79 DLH_X1 $T=55150 54200 0 0 $X=55035 $Y=54085
X3110 54 50 71 34 79 DLH_X1 $T=56100 59800 1 0 $X=55985 $Y=58285
X3111 67 79 56 62 61 114 34 NOR4_X1 $T=49260 59800 0 180 $X=48195 $Y=58285
X3112 64 79 252 254 71 138 34 NOR4_X1 $T=54390 57000 1 0 $X=54275 $Y=55485
X3113 63 196 60 201 68 34 79 NOR4_X2 $T=43180 59800 1 0 $X=43065 $Y=58285
X3136 81 2 156 263 34 79 AOI21_X1 $T=4610 54200 1 0 $X=4495 $Y=52685
X3137 301 9 266 325 34 79 AOI21_X1 $T=11830 54200 0 0 $X=11715 $Y=54085
X3138 268 23 303 265 34 79 AOI21_X1 $T=15820 54200 0 180 $X=14945 $Y=52685
X3139 98 107 187 212 34 79 AOI21_X1 $T=18670 51400 0 0 $X=18555 $Y=51285
X3140 93 29 270 309 34 79 AOI21_X1 $T=21140 51400 0 0 $X=21025 $Y=51285
X3141 327 27 341 180 34 79 AOI21_X1 $T=21900 54200 1 180 $X=21025 $Y=54085
X3142 221 27 328 331 34 79 AOI21_X1 $T=23040 57000 0 0 $X=22925 $Y=56885
X3143 98 32 279 167 34 79 AOI21_X1 $T=23990 59800 0 180 $X=23115 $Y=58285
X3144 98 36 278 181 34 79 AOI21_X1 $T=24750 59800 0 180 $X=23875 $Y=58285
X3145 222 27 343 311 34 79 AOI21_X1 $T=24750 57000 0 0 $X=24635 $Y=56885
X3146 98 19 313 158 34 79 AOI21_X1 $T=24750 59800 1 0 $X=24635 $Y=58285
X3147 55 228 280 344 34 79 AOI21_X1 $T=32730 57000 0 180 $X=31855 $Y=55485
X3148 349 246 168 345 34 79 AOI21_X1 $T=45840 54200 0 180 $X=44965 $Y=52685
X3149 247 248 349 292 34 79 AOI21_X1 $T=45840 54200 1 0 $X=45725 $Y=52685
X3152 149 6 34 213 264 79 85 212 OAI221_X1 $T=9740 51400 0 0 $X=9625 $Y=51285
X3153 86 6 34 214 7 79 11 265 OAI221_X1 $T=11450 59800 1 0 $X=11335 $Y=58285
X3154 127 85 34 216 217 79 6 87 OAI221_X1 $T=11830 51400 0 0 $X=11715 $Y=51285
X3155 220 29 34 26 31 79 28 329 OAI221_X1 $T=22280 54200 0 0 $X=22165 $Y=54085
X3156 229 280 34 230 231 79 11 242 OAI221_X1 $T=34060 57000 0 0 $X=33945 $Y=56885
X3157 156 1 79 122 298 123 34 AOI22_X1 $T=1950 54200 0 0 $X=1835 $Y=54085
X3158 299 1 79 122 347 34 34 AOI22_X1 $T=3280 57000 0 180 $X=2215 $Y=55485
X3159 298 146 79 172 217 145 34 AOI22_X1 $T=4610 54200 0 180 $X=3545 $Y=52685
X3160 298 172 79 146 147 121 34 AOI22_X1 $T=4040 51400 0 0 $X=3925 $Y=51285
X3161 262 3 79 82 173 148 34 AOI22_X1 $T=4990 59800 1 0 $X=4875 $Y=58285
X3162 15 20 79 92 124 17 34 AOI22_X1 $T=8600 54200 1 180 $X=7535 $Y=54085
X3163 15 25 79 88 262 17 34 AOI22_X1 $T=8030 57000 0 0 $X=7915 $Y=56885
X3164 15 12 79 78 80 17 34 AOI22_X1 $T=8220 57000 1 0 $X=8105 $Y=55485
X3165 15 18 79 91 148 17 34 AOI22_X1 $T=8980 57000 0 0 $X=8865 $Y=56885
X3166 264 9 79 125 213 149 34 AOI22_X1 $T=10120 54200 0 180 $X=9055 $Y=52685
X3167 15 13 79 16 174 17 34 AOI22_X1 $T=9550 59800 1 0 $X=9435 $Y=58285
X3168 86 125 79 11 214 98 34 AOI22_X1 $T=11450 59800 0 180 $X=10385 $Y=58285
X3169 127 9 79 125 216 217 34 AOI22_X1 $T=10880 51400 0 0 $X=10765 $Y=51285
X3170 126 125 79 8 215 98 34 AOI22_X1 $T=11640 57000 1 0 $X=11525 $Y=55485
X3171 267 150 79 129 301 302 34 AOI22_X1 $T=14110 54200 1 0 $X=13995 $Y=52685
X3172 267 129 79 150 264 128 34 AOI22_X1 $T=14490 51400 0 0 $X=14375 $Y=51285
X3173 271 129 79 150 22 302 34 AOI22_X1 $T=15820 54200 1 180 $X=14755 $Y=54085
X3174 270 27 79 26 271 304 34 AOI22_X1 $T=16770 54200 0 0 $X=16655 $Y=54085
X3175 271 150 79 129 199 326 34 AOI22_X1 $T=16960 59800 1 0 $X=16845 $Y=58285
X3176 269 129 79 150 175 219 34 AOI22_X1 $T=17530 57000 0 0 $X=17415 $Y=56885
X3177 304 27 79 26 219 305 34 AOI22_X1 $T=17720 54200 0 0 $X=17605 $Y=54085
X3178 306 129 79 150 218 269 34 AOI22_X1 $T=18670 57000 0 180 $X=17605 $Y=55485
X3179 219 129 79 150 177 326 34 AOI22_X1 $T=18860 59800 0 180 $X=17795 $Y=58285
X3180 176 27 79 26 302 340 34 AOI22_X1 $T=18100 54200 1 0 $X=17985 $Y=52685
X3181 328 129 79 150 178 306 34 AOI22_X1 $T=18480 57000 0 0 $X=18365 $Y=56885
X3182 305 27 79 26 306 273 34 AOI22_X1 $T=18670 57000 1 0 $X=18555 $Y=55485
X3183 340 27 79 26 326 276 34 AOI22_X1 $T=19430 54200 1 0 $X=19315 $Y=52685
X3184 179 29 79 28 307 312 34 AOI22_X1 $T=20380 54200 1 0 $X=20265 $Y=52685
X3185 273 27 79 26 275 327 34 AOI22_X1 $T=20950 57000 1 0 $X=20835 $Y=55485
X3186 275 129 79 150 94 328 34 AOI22_X1 $T=20950 59800 1 0 $X=20835 $Y=58285
X3187 275 150 79 129 131 308 34 AOI22_X1 $T=21140 57000 0 0 $X=21025 $Y=56885
X3188 341 329 79 150 157 308 34 AOI22_X1 $T=23040 57000 1 180 $X=21975 $Y=56885
X3189 276 27 79 26 269 221 34 AOI22_X1 $T=22280 57000 1 0 $X=22165 $Y=55485
X3190 31 28 79 29 353 312 34 AOI22_X1 $T=23420 54200 0 180 $X=22355 $Y=52685
X3191 96 28 79 29 310 133 34 AOI22_X1 $T=24180 51400 1 180 $X=23115 $Y=51285
X3192 330 29 79 28 277 33 34 AOI22_X1 $T=23420 54200 0 0 $X=23305 $Y=54085
X3193 224 28 79 29 342 97 34 AOI22_X1 $T=25320 54200 1 180 $X=24255 $Y=54085
X3194 97 28 79 29 354 34 34 AOI22_X1 $T=24940 54200 1 0 $X=24825 $Y=52685
X3195 159 28 79 29 222 96 34 AOI22_X1 $T=26460 51400 1 180 $X=25395 $Y=51285
X3196 38 103 79 41 312 99 34 AOI22_X1 $T=25890 54200 1 0 $X=25775 $Y=52685
X3197 38 35 79 49 34 99 34 AOI22_X1 $T=26460 51400 0 0 $X=26345 $Y=51285
X3198 38 40 79 225 330 99 34 AOI22_X1 $T=28550 51400 0 0 $X=28435 $Y=51285
X3199 104 227 79 283 281 223 34 AOI22_X1 $T=31780 54200 0 0 $X=31665 $Y=54085
X3200 281 315 79 42 344 282 34 AOI22_X1 $T=32730 54200 0 0 $X=32615 $Y=54085
X3201 106 19 79 48 289 134 34 AOI22_X1 $T=35010 51400 0 0 $X=34895 $Y=51285
X3202 106 39 79 226 232 134 34 AOI22_X1 $T=35010 54200 1 0 $X=34895 $Y=52685
X3203 50 235 79 233 230 48 34 AOI22_X1 $T=36150 57000 1 180 $X=35085 $Y=56885
X3204 106 21 79 55 287 134 34 AOI22_X1 $T=35960 51400 0 0 $X=35845 $Y=51285
X3205 251 333 79 288 245 290 34 AOI22_X1 $T=42420 54200 0 0 $X=42305 $Y=54085
X3206 113 59 79 161 248 137 34 AOI22_X1 $T=46030 51400 0 0 $X=45915 $Y=51285
X3207 301 85 34 325 6 126 79 OAI22_X1 $T=10880 54200 0 0 $X=10765 $Y=54085
X3208 44 234 34 229 228 55 79 OAI22_X1 $T=34060 57000 1 180 $X=32995 $Y=56885
X3209 288 290 34 291 334 243 79 OAI22_X1 $T=43180 57000 1 0 $X=43065 $Y=55485
X3210 251 333 34 316 317 318 79 OAI22_X1 $T=44320 54200 0 0 $X=44205 $Y=54085
X3222 348 28 79 27 33 34 29 311 AOI221_X1 $T=26460 57000 0 180 $X=25205 $Y=55485
X3223 225 284 79 236 49 34 188 109 AOI221_X1 $T=38810 51400 1 180 $X=37555 $Y=51285
X3224 241 8 79 237 239 34 36 236 AOI221_X1 $T=38430 54200 0 0 $X=38315 $Y=54085
X3225 285 32 79 240 238 34 10 332 AOI221_X1 $T=39760 57000 1 180 $X=38505 $Y=56885
X3226 34 1 145 261 34 79 34 OAI21_X1 $T=2330 59800 1 0 $X=2215 $Y=58285
X3227 262 3 299 324 34 79 34 OAI21_X1 $T=4800 57000 1 0 $X=4685 $Y=55485
X3228 124 3 34 300 34 79 34 OAI21_X1 $T=4800 57000 0 0 $X=4685 $Y=56885
X3229 268 24 251 303 34 79 34 OAI21_X1 $T=16200 51400 1 180 $X=15325 $Y=51285
X3230 270 27 267 272 34 79 34 OAI21_X1 $T=17340 51400 0 0 $X=17225 $Y=51285
X3231 130 28 340 274 34 79 34 OAI21_X1 $T=19430 51400 0 0 $X=19315 $Y=51285
X3232 7 10 288 195 34 79 34 OAI21_X1 $T=27600 59800 0 180 $X=26725 $Y=58285
X3233 7 36 160 278 34 79 34 OAI21_X1 $T=27980 57000 0 180 $X=27105 $Y=55485
X3234 7 19 317 313 34 79 34 OAI21_X1 $T=27220 57000 0 0 $X=27105 $Y=56885
X3235 7 32 334 279 34 79 34 OAI21_X1 $T=27600 59800 1 0 $X=27485 $Y=58285
X3236 7 39 101 100 34 79 34 OAI21_X1 $T=27980 57000 1 0 $X=27865 $Y=55485
X3237 7 42 113 102 34 79 34 OAI21_X1 $T=30450 57000 0 180 $X=29575 $Y=55485
X3238 7 21 161 152 34 79 34 OAI21_X1 $T=30450 57000 1 0 $X=30335 $Y=55485
X3239 46 226 58 232 34 79 34 OAI21_X1 $T=41090 51400 1 180 $X=40215 $Y=51285
X3240 46 55 137 287 34 79 34 OAI21_X1 $T=41090 51400 0 0 $X=40975 $Y=51285
X3241 46 48 318 289 34 79 34 OAI21_X1 $T=42230 54200 1 0 $X=42115 $Y=52685
X3242 291 245 345 319 34 79 34 OAI21_X1 $T=44130 57000 1 0 $X=44015 $Y=55485
X3243 34 34 1 261 79 NAND2_X1 $T=2330 57000 0 0 $X=2215 $Y=56885
X3244 81 34 18 324 79 NAND2_X1 $T=6130 57000 0 180 $X=5445 $Y=55485
X3245 81 34 83 300 79 NAND2_X1 $T=6700 57000 0 0 $X=6585 $Y=56885
X3246 186 34 27 272 79 NAND2_X1 $T=18670 51400 1 180 $X=17985 $Y=51285
X3247 330 34 28 274 79 NAND2_X1 $T=23990 54200 0 180 $X=23305 $Y=52685
X3248 243 34 334 319 79 NAND2_X1 $T=45460 57000 0 180 $X=44775 $Y=55485
X3249 299 79 1 144 34 NOR2_X1 $T=2900 51400 1 180 $X=2215 $Y=51285
X3250 80 79 3 263 34 NOR2_X1 $T=6130 54200 1 180 $X=5445 $Y=54085
X3251 5 79 4 14 34 NOR2_X1 $T=12590 54200 0 0 $X=12475 $Y=54085
X3252 34 79 29 309 34 NOR2_X1 $T=22280 51400 0 0 $X=22165 $Y=51285
X3253 222 79 27 331 34 NOR2_X1 $T=24750 57000 1 180 $X=24065 $Y=56885
X3254 316 79 291 246 34 NOR2_X1 $T=44510 54200 1 0 $X=44395 $Y=52685
X3255 137 79 161 292 34 NOR2_X1 $T=47550 51400 1 180 $X=46865 $Y=51285
X3256 57 79 66 253 34 154 NOR3_X1 $T=51730 51400 0 0 $X=51615 $Y=51285
X3259 350 293 318 317 79 34 153 FA_X1 $T=48310 54200 1 180 $X=45155 $Y=54085
X3260 249 350 290 288 79 34 115 FA_X1 $T=45460 57000 1 0 $X=45345 $Y=55485
X3261 293 251 333 349 79 34 117 FA_X1 $T=47550 51400 0 0 $X=47435 $Y=51285
X3262 34 243 250 249 79 XNOR2_X1 $T=46030 57000 0 0 $X=45915 $Y=56885
X3263 34 334 197 250 79 XNOR2_X1 $T=48310 57000 1 180 $X=47055 $Y=56885
X3265 7 8 266 79 215 200 34 OAI211_X1 $T=12780 54200 0 180 $X=11715 $Y=52685
X3266 7 30 132 79 95 151 34 OAI211_X1 $T=23230 59800 0 180 $X=22165 $Y=58285
X3267 104 227 314 79 226 315 34 OAI211_X1 $T=31780 54200 1 0 $X=31665 $Y=52685
X3268 113 59 101 79 58 247 34 OAI211_X1 $T=45080 51400 1 180 $X=44015 $Y=51285
X3269 108 282 34 223 46 47 79 283 59 OAI222_X1 $T=34820 54200 0 0 $X=34705 $Y=54085
X3270 108 231 34 44 46 47 79 234 333 OAI222_X1 $T=35770 57000 1 0 $X=35655 $Y=55485
X3271 108 238 34 50 46 47 79 235 290 OAI222_X1 $T=38810 57000 0 180 $X=37175 $Y=55485
X3272 108 241 34 225 46 47 79 284 135 OAI222_X1 $T=38810 51400 0 0 $X=38695 $Y=51285
X3273 108 239 34 41 46 47 79 244 136 OAI222_X1 $T=39950 54200 0 0 $X=39835 $Y=54085
X3274 108 285 34 51 46 47 79 286 243 OAI222_X1 $T=40330 57000 1 0 $X=40215 $Y=55485
X3275 50 235 48 34 233 240 79 AOI211_X1 $T=37100 57000 1 180 $X=36035 $Y=56885
X3279 4 17 84 34 79 NOR2_X2 $T=9170 54200 0 180 $X=8105 $Y=52685
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 A3 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI33_X1 B3 B2 B1 VSS A1 A2 A3 ZN VDD
** N=14 EP=9 IP=0 FDC=12
M0 10 B3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS B2 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 10 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 10 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 ZN A3 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1110 $Y=90 $D=1
M6 11 B3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M7 12 B2 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M8 ZN B1 12 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M9 13 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M10 14 A2 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
M11 VDD A3 14 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1110 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221
+ 222
** N=367 EP=221 IP=5312 FDC=2024
X2624 186 50 85 86 44 85 DFF_X1 $T=42230 43000 1 0 $X=42115 $Y=41485
X2625 343 73 85 86 61 85 DFF_X1 $T=58760 51400 1 0 $X=58645 $Y=49885
X2626 324 83 85 86 171 85 DFF_X1 $T=65790 43000 1 0 $X=65675 $Y=41485
X2627 357 73 85 86 47 85 DFF_X1 $T=65790 45800 1 0 $X=65675 $Y=44285
X2628 355 73 85 86 119 85 DFF_X1 $T=65790 48600 1 0 $X=65675 $Y=47085
X2629 296 83 85 86 180 85 DFF_X1 $T=66170 45800 0 0 $X=66055 $Y=45685
X2630 187 83 85 86 172 85 DFF_X1 $T=66170 51400 1 0 $X=66055 $Y=49885
X2709 128 62 85 86 296 85 AND2_X1 $T=51160 45800 1 0 $X=51045 $Y=44285
X2710 169 65 85 86 126 85 AND2_X1 $T=53820 51400 1 0 $X=53705 $Y=49885
X2711 170 74 85 86 262 85 AND2_X1 $T=60470 43000 1 0 $X=60355 $Y=41485
X2712 128 263 85 86 324 85 AND2_X1 $T=61230 43000 1 0 $X=61115 $Y=41485
X2713 129 80 85 86 355 85 AND2_X1 $T=64270 45800 0 0 $X=64155 $Y=45685
X2714 129 81 85 86 343 85 AND2_X1 $T=64270 51400 1 0 $X=64155 $Y=49885
X2715 129 82 85 86 357 85 AND2_X1 $T=65030 43000 1 0 $X=64915 $Y=41485
X3186 270 85 86 269 85 INV_X1 $T=8030 43000 1 0 $X=7915 $Y=41485
X3187 268 85 86 358 85 INV_X1 $T=8030 43000 0 0 $X=7915 $Y=42885
X3188 204 85 86 3 85 INV_X1 $T=8790 51400 0 180 $X=8295 $Y=49885
X3189 134 85 86 5 85 INV_X1 $T=9360 43000 0 0 $X=9245 $Y=42885
X3190 4 85 86 133 85 INV_X1 $T=9360 51400 1 0 $X=9245 $Y=49885
X3191 136 85 86 9 85 INV_X1 $T=13540 43000 1 180 $X=13045 $Y=42885
X3192 7 85 86 97 85 INV_X1 $T=13540 43000 0 0 $X=13425 $Y=42885
X3193 153 85 86 96 85 INV_X1 $T=16010 51400 0 180 $X=15515 $Y=49885
X3194 104 85 86 18 85 INV_X1 $T=22280 43000 0 0 $X=22165 $Y=42885
X3195 16 85 86 17 85 INV_X1 $T=22660 48600 1 180 $X=22165 $Y=48485
X3196 92 85 86 238 85 INV_X1 $T=22660 43000 0 0 $X=22545 $Y=42885
X3197 159 85 86 313 85 INV_X1 $T=23990 45800 0 180 $X=23495 $Y=44285
X3198 22 85 86 287 85 INV_X1 $T=23610 45800 0 0 $X=23495 $Y=45685
X3199 102 85 86 23 85 INV_X1 $T=24370 45800 1 0 $X=24255 $Y=44285
X3200 25 85 86 240 85 INV_X1 $T=25130 43000 1 0 $X=25015 $Y=41485
X3201 35 85 86 242 85 INV_X1 $T=27600 43000 0 0 $X=27485 $Y=42885
X3202 24 85 86 332 85 INV_X1 $T=27790 48600 1 0 $X=27675 $Y=47085
X3203 31 85 86 246 85 INV_X1 $T=29120 43000 1 0 $X=29005 $Y=41485
X3204 36 85 86 333 85 INV_X1 $T=30450 48600 0 180 $X=29955 $Y=47085
X3205 15 85 86 247 85 INV_X1 $T=30640 43000 1 180 $X=30145 $Y=42885
X3206 42 85 86 245 85 INV_X1 $T=31210 45800 1 180 $X=30715 $Y=45685
X3207 43 85 86 291 85 INV_X1 $T=31780 48600 0 0 $X=31665 $Y=48485
X3208 12 85 86 248 85 INV_X1 $T=32920 48600 0 180 $X=32425 $Y=47085
X3209 45 85 86 113 85 INV_X1 $T=32920 48600 0 0 $X=32805 $Y=48485
X3210 14 85 86 292 85 INV_X1 $T=35390 48600 0 180 $X=34895 $Y=47085
X3211 115 85 86 212 85 INV_X1 $T=35200 45800 0 0 $X=35085 $Y=45685
X3212 243 85 86 318 85 INV_X1 $T=35390 48600 1 0 $X=35275 $Y=47085
X3213 116 85 86 319 85 INV_X1 $T=35960 51400 0 180 $X=35465 $Y=49885
X3214 207 85 86 118 85 INV_X1 $T=37290 45800 0 0 $X=37175 $Y=45685
X3215 143 85 86 362 85 INV_X1 $T=38050 48600 1 180 $X=37555 $Y=48485
X3216 39 85 86 144 85 INV_X1 $T=38050 48600 0 0 $X=37935 $Y=48485
X3217 208 85 86 85 85 INV_X1 $T=39000 51400 1 0 $X=38885 $Y=49885
X3218 347 85 86 353 85 INV_X1 $T=40330 45800 1 0 $X=40215 $Y=44285
X3219 119 85 86 145 85 INV_X1 $T=43560 45800 0 0 $X=43445 $Y=45685
X3220 209 85 86 349 85 INV_X1 $T=44890 51400 0 180 $X=44395 $Y=49885
X3221 356 85 86 148 85 INV_X1 $T=50020 48600 0 0 $X=49905 $Y=48485
X3222 366 85 86 185 85 INV_X1 $T=50780 48600 0 0 $X=50665 $Y=48485
X3223 341 85 86 263 85 INV_X1 $T=53060 43000 1 0 $X=52945 $Y=41485
X3224 302 85 86 350 85 INV_X1 $T=58190 51400 0 180 $X=57695 $Y=49885
X3333 205 238 86 9 239 8 85 92 367 AOI222_X1 $T=19430 43000 0 0 $X=19315 $Y=42885
X3334 38 108 86 19 20 21 85 43 109 AOI222_X1 $T=22660 48600 0 0 $X=22545 $Y=48485
X3335 38 26 86 28 20 21 85 35 110 AOI222_X1 $T=25700 48600 1 0 $X=25585 $Y=47085
X3336 38 215 86 32 20 21 85 243 175 AOI222_X1 $T=26840 51400 1 0 $X=26725 $Y=49885
X3337 38 33 86 34 20 21 85 42 206 AOI222_X1 $T=27790 48600 0 0 $X=27675 $Y=48485
X3338 21 36 86 37 38 20 85 107 184 AOI222_X1 $T=28360 51400 1 0 $X=28245 $Y=49885
X3339 51 47 86 53 44 54 85 178 341 AOI222_X1 $T=45460 43000 1 0 $X=45345 $Y=41485
X3340 120 59 86 58 57 56 85 121 356 AOI222_X1 $T=50400 45800 1 180 $X=48765 $Y=45685
X3341 120 58 86 60 57 56 85 295 366 AOI222_X1 $T=49450 43000 0 0 $X=49335 $Y=42885
X3342 120 258 86 59 57 56 85 297 124 AOI222_X1 $T=50590 48600 1 0 $X=50475 $Y=47085
X3343 120 261 86 260 57 56 85 298 125 AOI222_X1 $T=55150 45800 1 180 $X=53515 $Y=45685
X3344 120 64 86 258 57 56 85 299 211 AOI222_X1 $T=55150 48600 1 180 $X=53515 $Y=48485
X3345 120 260 86 67 57 56 85 365 127 AOI222_X1 $T=55150 45800 0 0 $X=55035 $Y=45685
X3346 120 63 86 64 57 56 85 325 202 AOI222_X1 $T=55150 48600 0 0 $X=55035 $Y=48485
X3347 51 61 86 53 71 54 85 350 216 AOI222_X1 $T=56290 51400 1 0 $X=56175 $Y=49885
X3348 120 69 86 261 57 56 85 300 302 AOI222_X1 $T=56670 45800 0 0 $X=56555 $Y=45685
X3349 120 70 86 63 57 56 85 301 217 AOI222_X1 $T=56670 48600 0 0 $X=56555 $Y=48485
X3350 120 67 86 70 57 56 85 342 218 AOI222_X1 $T=57430 48600 1 0 $X=57315 $Y=47085
X3375 195 12 40 85 86 DLH_X1 $T=29500 43000 1 0 $X=29385 $Y=41485
X3376 54 14 44 85 86 DLH_X1 $T=31780 45800 1 0 $X=31665 $Y=44285
X3377 54 198 46 85 86 DLH_X1 $T=34630 51400 0 180 $X=32615 $Y=49885
X3378 54 243 47 85 86 DLH_X1 $T=37290 45800 1 0 $X=37175 $Y=44285
X3379 56 123 258 85 86 DLH_X1 $T=49450 43000 1 180 $X=47435 $Y=42885
X3380 54 48 61 85 86 DLH_X1 $T=50210 51400 1 0 $X=50095 $Y=49885
X3381 56 85 63 85 86 DLH_X1 $T=50400 45800 0 0 $X=50285 $Y=45685
X3382 56 170 259 85 86 DLH_X1 $T=51160 43000 1 0 $X=51045 $Y=41485
X3383 56 179 64 85 86 DLH_X1 $T=51920 43000 0 0 $X=51805 $Y=42885
X3384 56 220 260 85 86 DLH_X1 $T=53630 45800 1 0 $X=53515 $Y=44285
X3385 149 298 66 85 86 DLH_X1 $T=56290 43000 0 180 $X=54275 $Y=41485
X3386 149 365 68 85 86 DLH_X1 $T=56100 43000 0 0 $X=55985 $Y=42885
X3387 56 203 261 85 86 DLH_X1 $T=58570 43000 1 0 $X=58455 $Y=41485
X3388 149 301 72 85 86 DLH_X1 $T=58950 48600 1 0 $X=58835 $Y=47085
X3389 149 300 262 85 86 DLH_X1 $T=61990 43000 1 180 $X=59975 $Y=42885
X3390 149 342 75 85 86 DLH_X1 $T=61990 45800 1 180 $X=59975 $Y=45685
X3391 56 150 70 85 86 DLH_X1 $T=60090 48600 0 0 $X=59975 $Y=48485
X3392 149 295 76 85 86 DLH_X1 $T=61990 43000 0 0 $X=61875 $Y=42885
X3393 149 297 77 85 86 DLH_X1 $T=62370 45800 1 0 $X=62255 $Y=44285
X3394 149 299 78 85 86 DLH_X1 $T=62370 45800 0 0 $X=62255 $Y=45685
X3395 149 325 79 85 86 DLH_X1 $T=62370 48600 0 0 $X=62255 $Y=48485
X3396 46 86 161 71 163 162 85 NOR4_X1 $T=31400 43000 1 0 $X=31285 $Y=41485
X3413 305 1 264 181 85 86 AOI21_X1 $T=1190 48600 0 0 $X=1075 $Y=48485
X3414 307 9 308 306 85 86 AOI21_X1 $T=11450 43000 0 0 $X=11335 $Y=42885
X3415 8 12 331 326 85 86 AOI21_X1 $T=16960 48600 0 180 $X=16085 $Y=47085
X3416 328 13 275 281 85 86 AOI21_X1 $T=16200 48600 0 0 $X=16085 $Y=48485
X3417 8 24 288 359 85 86 AOI21_X1 $T=16770 45800 0 0 $X=16655 $Y=45685
X3418 8 15 289 284 85 86 AOI21_X1 $T=16960 48600 1 0 $X=16845 $Y=47085
X3419 8 14 290 194 85 86 AOI21_X1 $T=17720 51400 0 180 $X=16845 $Y=49885
X3420 103 18 241 351 85 86 AOI21_X1 $T=23800 43000 0 0 $X=23685 $Y=42885
X3421 23 10 351 352 85 86 AOI21_X1 $T=24560 43000 0 0 $X=24445 $Y=42885
X3422 43 248 244 344 85 86 AOI21_X1 $T=31780 48600 1 0 $X=31665 $Y=47085
X3423 291 12 344 335 85 86 AOI21_X1 $T=32160 48600 0 0 $X=32045 $Y=48485
X3424 353 250 176 345 85 86 AOI21_X1 $T=37860 43000 1 180 $X=36985 $Y=42885
X3425 349 253 347 339 85 86 AOI21_X1 $T=40710 48600 0 180 $X=39835 $Y=47085
X3429 227 7 85 228 229 86 5 359 OAI221_X1 $T=9170 45800 0 0 $X=9055 $Y=45685
X3430 267 5 85 230 231 86 7 284 OAI221_X1 $T=9740 48600 1 0 $X=9625 $Y=47085
X3431 272 7 85 233 6 86 5 326 OAI221_X1 $T=11260 48600 1 180 $X=10005 $Y=48485
X3432 273 7 85 234 232 86 5 235 OAI221_X1 $T=11450 45800 1 180 $X=10195 $Y=45685
X3433 23 10 85 241 240 86 92 222 OAI221_X1 $T=24370 43000 0 180 $X=23115 $Y=41485
X3434 245 15 85 244 242 86 31 361 OAI221_X1 $T=29310 45800 0 180 $X=28055 $Y=44285
X3435 264 133 86 87 229 304 85 AOI22_X1 $T=2140 45800 0 0 $X=2025 $Y=45685
X3436 188 1 86 131 266 305 85 AOI22_X1 $T=2330 43000 0 0 $X=2215 $Y=42885
X3437 189 1 86 131 304 265 85 AOI22_X1 $T=2330 45800 1 0 $X=2215 $Y=44285
X3438 304 133 86 87 271 266 85 AOI22_X1 $T=3280 43000 0 0 $X=3165 $Y=42885
X3439 264 87 86 133 232 303 85 AOI22_X1 $T=3660 48600 0 0 $X=3545 $Y=48485
X3440 88 132 86 10 265 91 85 AOI22_X1 $T=4610 48600 0 0 $X=4495 $Y=48485
X3441 88 90 86 104 189 91 85 AOI22_X1 $T=4800 45800 0 0 $X=4685 $Y=45685
X3442 182 133 86 221 270 87 85 AOI22_X1 $T=5180 43000 1 0 $X=5065 $Y=41485
X3443 89 133 86 87 267 303 85 AOI22_X1 $T=5370 51400 1 0 $X=5255 $Y=49885
X3444 182 87 86 133 268 266 85 AOI22_X1 $T=5750 43000 0 0 $X=5635 $Y=42885
X3445 91 84 86 190 188 88 85 AOI22_X1 $T=6510 45800 1 0 $X=6395 $Y=44285
X3446 88 93 86 92 305 91 85 AOI22_X1 $T=7080 48600 1 0 $X=6965 $Y=47085
X3447 229 135 86 9 228 227 85 AOI22_X1 $T=8220 45800 0 0 $X=8105 $Y=45685
X3448 269 134 86 135 191 270 85 AOI22_X1 $T=8410 43000 1 0 $X=8295 $Y=41485
X3449 358 134 86 135 237 268 85 AOI22_X1 $T=9360 43000 1 180 $X=8295 $Y=42885
X3450 267 135 86 9 230 231 85 AOI22_X1 $T=9170 48600 0 0 $X=9055 $Y=48485
X3451 272 9 86 135 233 6 85 AOI22_X1 $T=9740 51400 1 0 $X=9625 $Y=49885
X3452 271 135 86 10 236 8 85 AOI22_X1 $T=10690 43000 1 0 $X=10575 $Y=41485
X3453 276 96 86 152 273 274 85 AOI22_X1 $T=13350 48600 0 180 $X=12285 $Y=47085
X3454 275 96 86 152 272 277 85 AOI22_X1 $T=12780 48600 0 0 $X=12665 $Y=48485
X3455 276 152 86 96 231 277 85 AOI22_X1 $T=13350 48600 1 0 $X=13235 $Y=47085
X3456 275 152 86 96 137 98 85 AOI22_X1 $T=13350 51400 1 0 $X=13235 $Y=49885
X3457 274 96 86 152 227 309 85 AOI22_X1 $T=13540 45800 0 0 $X=13425 $Y=45685
X3458 13 28 86 19 193 99 85 AOI22_X1 $T=13920 43000 1 0 $X=13805 $Y=41485
X3459 309 96 86 152 307 310 85 AOI22_X1 $T=13920 45800 1 0 $X=13805 $Y=44285
X3460 279 13 86 99 274 327 85 AOI22_X1 $T=14300 48600 1 0 $X=14185 $Y=47085
X3461 282 13 86 99 309 311 85 AOI22_X1 $T=14490 45800 0 0 $X=14375 $Y=45685
X3462 278 13 86 99 310 279 85 AOI22_X1 $T=14870 45800 1 0 $X=14755 $Y=44285
X3463 311 13 86 99 276 328 85 AOI22_X1 $T=15250 48600 1 0 $X=15135 $Y=47085
X3464 327 13 86 99 277 312 85 AOI22_X1 $T=15250 48600 0 0 $X=15135 $Y=48485
X3465 312 13 86 99 98 11 85 AOI22_X1 $T=16960 51400 0 180 $X=15895 $Y=49885
X3466 152 138 86 96 183 283 85 AOI22_X1 $T=16390 43000 1 0 $X=16275 $Y=41485
X3467 286 107 86 32 278 100 85 AOI22_X1 $T=18480 45800 0 180 $X=17415 $Y=44285
X3468 286 34 86 25 279 100 85 AOI22_X1 $T=18480 45800 1 180 $X=17415 $Y=45685
X3469 152 283 86 96 239 310 85 AOI22_X1 $T=18480 43000 0 0 $X=18365 $Y=42885
X3470 286 28 86 103 282 100 85 AOI22_X1 $T=19430 45800 0 180 $X=18365 $Y=44285
X3471 286 32 86 17 327 285 85 AOI22_X1 $T=19810 48600 0 180 $X=18745 $Y=47085
X3472 286 19 86 102 311 100 85 AOI22_X1 $T=19620 45800 0 0 $X=19505 $Y=45685
X3473 286 25 86 17 312 140 85 AOI22_X1 $T=19620 48600 0 0 $X=19505 $Y=48485
X3474 286 103 86 17 328 157 85 AOI22_X1 $T=19810 48600 1 0 $X=19695 $Y=47085
X3475 21 19 86 43 155 38 85 AOI22_X1 $T=24180 48600 0 0 $X=24065 $Y=48485
X3476 21 32 86 243 158 38 85 AOI22_X1 $T=26840 48600 0 0 $X=26725 $Y=48485
X3477 360 361 86 332 352 36 85 AOI22_X1 $T=28360 45800 0 0 $X=28245 $Y=45685
X3478 197 196 86 48 340 112 85 AOI22_X1 $T=32730 51400 0 180 $X=31665 $Y=49885
X3479 251 316 86 30 249 142 85 AOI22_X1 $T=35390 43000 1 180 $X=34325 $Y=42885
X3480 243 292 86 362 335 317 85 AOI22_X1 $T=35580 48600 1 180 $X=34515 $Y=48485
X3481 319 39 86 14 317 318 85 AOI22_X1 $T=34630 51400 1 0 $X=34515 $Y=49885
X3482 49 199 86 338 252 322 85 AOI22_X1 $T=40710 48600 1 180 $X=39645 $Y=48485
X3483 57 69 86 259 201 120 85 AOI22_X1 $T=46980 43000 1 0 $X=46865 $Y=41485
X3484 265 131 85 303 1 151 86 OAI22_X1 $T=1950 51400 1 0 $X=1835 $Y=49885
X3485 307 7 85 306 5 271 86 OAI22_X1 $T=11450 43000 1 180 $X=10385 $Y=42885
X3486 278 13 85 138 139 280 86 OAI22_X1 $T=14870 43000 0 0 $X=14755 $Y=42885
X3487 280 154 85 283 13 282 86 OAI22_X1 $T=17530 43000 0 0 $X=17415 $Y=42885
X3488 30 142 85 334 164 114 86 OAI22_X1 $T=33490 43000 1 0 $X=33375 $Y=41485
X3489 251 316 85 293 141 41 86 OAI22_X1 $T=38810 43000 1 180 $X=37745 $Y=42885
X3490 338 322 85 294 323 321 86 OAI22_X1 $T=39190 48600 0 180 $X=38125 $Y=47085
X3491 49 199 85 320 166 165 86 OAI22_X1 $T=40330 51400 0 180 $X=39265 $Y=49885
X3495 232 135 86 235 8 85 31 314 AOI221_X1 $T=11070 45800 1 0 $X=10955 $Y=44285
X3496 333 24 86 315 242 85 31 360 AOI221_X1 $T=27030 45800 1 0 $X=26915 $Y=44285
X3497 155 16 101 329 85 86 85 OAI21_X1 $T=20380 51400 1 0 $X=20265 $Y=49885
X3498 285 17 11 330 85 86 85 OAI21_X1 $T=21140 51400 1 0 $X=21025 $Y=49885
X3499 117 23 160 173 85 86 85 OAI21_X1 $T=24370 43000 1 0 $X=24255 $Y=41485
X3500 95 12 251 331 85 86 85 OAI21_X1 $T=25700 48600 0 180 $X=24825 $Y=47085
X3501 95 24 164 288 85 86 85 OAI21_X1 $T=26270 45800 1 180 $X=25395 $Y=45685
X3502 95 15 141 289 85 86 85 OAI21_X1 $T=26270 45800 1 0 $X=26155 $Y=44285
X3503 95 31 30 314 85 86 85 OAI21_X1 $T=26840 43000 0 0 $X=26725 $Y=42885
X3504 95 39 338 111 85 86 85 OAI21_X1 $T=29880 51400 1 0 $X=29765 $Y=49885
X3505 95 14 323 290 85 86 85 OAI21_X1 $T=30070 48600 0 0 $X=29955 $Y=48485
X3506 334 249 345 336 85 86 85 OAI21_X1 $T=36530 43000 0 180 $X=35655 $Y=41485
X3507 294 252 339 337 85 86 85 OAI21_X1 $T=39190 48600 1 0 $X=39075 $Y=47085
X3508 27 48 364 340 85 86 85 OAI21_X1 $T=41850 51400 1 0 $X=41735 $Y=49885
X3509 273 85 9 234 86 NAND2_X1 $T=11450 48600 0 180 $X=10765 $Y=47085
X3510 13 85 100 280 86 NAND2_X1 $T=15820 43000 0 0 $X=15705 $Y=42885
X3511 286 85 102 329 86 NAND2_X1 $T=20570 48600 0 0 $X=20455 $Y=48485
X3512 158 85 17 330 86 NAND2_X1 $T=23420 51400 0 180 $X=22735 $Y=49885
X3513 114 85 164 336 86 NAND2_X1 $T=35200 43000 1 0 $X=35085 $Y=41485
X3514 321 85 323 337 86 NAND2_X1 $T=37670 48600 1 0 $X=37555 $Y=47085
X3515 101 86 13 281 85 NOR2_X1 $T=18290 51400 0 180 $X=17605 $Y=49885
X3516 313 86 287 21 85 NOR2_X1 $T=24370 48600 0 180 $X=23685 $Y=47085
X3517 159 86 22 20 85 NOR2_X1 $T=24560 45800 1 180 $X=23875 $Y=45685
X3518 313 86 22 38 85 NOR2_X1 $T=24370 48600 1 0 $X=24255 $Y=47085
X3519 293 86 334 250 85 NOR2_X1 $T=37100 43000 0 180 $X=36415 $Y=41485
X3520 320 86 294 253 85 NOR2_X1 $T=39000 48600 1 180 $X=38315 $Y=48485
X3521 94 86 3 2 85 91 NOR3_X1 $T=8410 51400 0 180 $X=7535 $Y=49885
X3522 17 86 313 22 85 286 NOR3_X1 $T=20760 48600 1 0 $X=20645 $Y=47085
X3523 16 86 313 22 85 100 NOR3_X1 $T=21710 43000 1 180 $X=20835 $Y=42885
X3525 177 251 316 353 86 85 200 FA_X1 $T=38810 43000 0 0 $X=38695 $Y=42885
X3526 346 363 322 338 86 85 58 FA_X1 $T=39570 45800 0 0 $X=39455 $Y=45685
X3527 363 348 165 166 86 85 59 FA_X1 $T=42230 48600 1 0 $X=42115 $Y=47085
X3528 348 49 199 349 86 85 258 FA_X1 $T=42230 48600 0 0 $X=42115 $Y=48485
X3529 255 52 219 85 86 85 259 FA_X1 $T=46410 45800 0 180 $X=43255 $Y=44285
X3530 256 255 364 213 86 85 69 FA_X1 $T=46980 45800 1 180 $X=43825 $Y=45685
X3531 257 256 214 210 86 85 261 FA_X1 $T=48310 48600 0 180 $X=45155 $Y=47085
X3532 85 321 254 346 86 XNOR2_X1 $T=39190 45800 1 0 $X=39075 $Y=44285
X3533 85 323 60 254 86 XNOR2_X1 $T=43370 45800 0 180 $X=42115 $Y=44285
X3534 85 167 354 257 86 XNOR2_X1 $T=46600 48600 0 0 $X=46485 $Y=48485
X3535 85 55 260 354 86 XNOR2_X1 $T=49260 51400 0 180 $X=48005 $Y=49885
X3538 95 10 308 86 236 192 85 OAI211_X1 $T=12590 43000 0 180 $X=11525 $Y=41485
X3539 239 7 237 86 367 86 85 OAI211_X1 $T=19240 43000 1 0 $X=19125 $Y=41485
X3540 117 240 85 25 27 29 86 238 174 OAI222_X1 $T=25510 43000 1 0 $X=25395 $Y=41485
X3541 117 242 85 35 27 29 86 246 142 OAI222_X1 $T=27980 43000 0 0 $X=27865 $Y=42885
X3542 117 333 85 36 27 29 86 332 114 OAI222_X1 $T=30830 45800 1 180 $X=29195 $Y=45685
X3543 117 245 85 42 27 29 86 247 41 OAI222_X1 $T=30260 45800 1 0 $X=30145 $Y=44285
X3544 117 291 85 43 27 29 86 248 316 OAI222_X1 $T=31210 45800 0 0 $X=31095 $Y=45685
X3545 117 318 85 243 27 29 86 292 321 OAI222_X1 $T=37670 48600 0 180 $X=36035 $Y=47085
X3546 117 319 85 116 27 29 86 144 322 OAI222_X1 $T=37480 51400 1 0 $X=37365 $Y=49885
X3547 103 18 25 85 238 106 86 AOI211_X1 $T=22280 43000 1 0 $X=22165 $Y=41485
X3548 35 246 42 85 247 315 86 AOI211_X1 $T=29310 45800 1 0 $X=29195 $Y=44285
X3555 168 85 146 147 122 86 86 NAND4_X1 $T=49260 51400 1 0 $X=49145 $Y=49885
X3558 156 313 287 85 22 313 242 157 86 OAI33_X1 $T=20570 45800 1 0 $X=20455 $Y=44285
X3559 139 313 287 85 22 313 245 140 86 OAI33_X1 $T=20570 45800 0 0 $X=20455 $Y=45685
X3560 105 313 287 85 22 313 333 285 86 OAI33_X1 $T=22280 45800 1 0 $X=22165 $Y=44285
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT BUF_X2 A Z VSS VDD
** N=5 EP=4 IP=0 FDC=6
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 5 Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VDD A 5 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD 5 Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X3 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=8
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 5 Z VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=715 $Y=90 $D=1
M4 VDD A 5 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 VDD 5 Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224
** N=357 EP=222 IP=4852 FDC=1840
X2345 350 2 101 71 7 101 DFF_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X2346 3 4 101 71 148 101 DFF_X1 $T=2330 34600 1 0 $X=2215 $Y=33085
X2347 351 2 101 71 6 101 DFF_X1 $T=2330 37400 0 0 $X=2215 $Y=37285
X2348 323 4 101 71 259 101 DFF_X1 $T=27600 34600 1 0 $X=27485 $Y=33085
X2417 102 182 101 71 322 101 AND2_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X2418 102 1 101 71 352 101 AND2_X1 $T=1190 34600 1 0 $X=1075 $Y=33085
X2419 147 5 101 71 323 101 AND2_X1 $T=3660 34600 0 0 $X=3545 $Y=34485
X2420 8 11 101 71 186 101 AND2_X1 $T=10120 40200 0 0 $X=10005 $Y=40085
X2421 8 14 101 71 105 101 AND2_X1 $T=12970 40200 0 0 $X=12855 $Y=40085
X2875 17 101 71 252 101 INV_X1 $T=6130 40200 0 180 $X=5635 $Y=38685
X2876 104 101 71 249 101 INV_X1 $T=7840 37400 1 180 $X=7345 $Y=37285
X2877 157 101 71 237 101 INV_X1 $T=11070 37400 1 0 $X=10955 $Y=35885
X2878 307 101 71 240 101 INV_X1 $T=11070 40200 0 0 $X=10955 $Y=40085
X2879 310 101 71 238 101 INV_X1 $T=12020 34600 0 0 $X=11905 $Y=34485
X2880 9 101 71 244 101 INV_X1 $T=15250 34600 1 180 $X=14755 $Y=34485
X2881 24 101 71 109 101 INV_X1 $T=17150 40200 0 0 $X=17035 $Y=40085
X2882 324 101 71 110 101 INV_X1 $T=18100 34600 1 0 $X=17985 $Y=33085
X2883 16 101 71 158 101 INV_X1 $T=18290 37400 1 0 $X=18175 $Y=35885
X2884 30 101 71 19 101 INV_X1 $T=18670 40200 0 180 $X=18175 $Y=38685
X2885 112 101 71 156 101 INV_X1 $T=19240 40200 0 0 $X=19125 $Y=40085
X2886 21 101 71 253 101 INV_X1 $T=20950 37400 0 0 $X=20835 $Y=37285
X2887 31 101 71 255 101 INV_X1 $T=21330 37400 0 0 $X=21215 $Y=37285
X2888 114 101 71 113 101 INV_X1 $T=22660 34600 0 180 $X=22165 $Y=33085
X2889 35 101 71 254 101 INV_X1 $T=23040 40200 1 180 $X=22545 $Y=40085
X2890 25 101 71 172 101 INV_X1 $T=23610 34600 1 180 $X=23115 $Y=34485
X2891 292 101 71 180 101 INV_X1 $T=27220 34600 1 0 $X=27105 $Y=33085
X2892 111 101 71 117 101 INV_X1 $T=30260 37400 0 0 $X=30145 $Y=37285
X2893 209 101 71 326 101 INV_X1 $T=32160 40200 1 0 $X=32045 $Y=38685
X2894 327 101 71 315 101 INV_X1 $T=36910 37400 0 180 $X=36415 $Y=35885
X2895 316 101 71 124 101 INV_X1 $T=37290 34600 0 0 $X=37175 $Y=34485
X2896 101 101 71 204 101 INV_X1 $T=40710 40200 1 0 $X=40595 $Y=38685
X2897 83 101 71 61 101 INV_X1 $T=42230 34600 0 0 $X=42115 $Y=34485
X2898 161 101 71 329 101 INV_X1 $T=43940 40200 1 180 $X=43445 $Y=40085
X2899 60 101 71 85 101 INV_X1 $T=46030 34600 1 0 $X=45915 $Y=33085
X2900 356 101 71 162 101 INV_X1 $T=46220 40200 0 0 $X=46105 $Y=40085
X2901 348 101 71 130 101 INV_X1 $T=49450 34600 1 0 $X=49335 $Y=33085
X2902 136 101 71 142 101 INV_X1 $T=58000 37400 1 0 $X=57885 $Y=35885
X2903 273 101 71 319 101 INV_X1 $T=58760 37400 0 180 $X=58265 $Y=35885
X2904 89 101 71 87 101 INV_X1 $T=60660 37400 0 0 $X=60545 $Y=37285
X2905 94 101 71 135 101 INV_X1 $T=64650 37400 0 180 $X=64155 $Y=35885
X2906 91 101 71 80 101 INV_X1 $T=65030 37400 0 180 $X=64535 $Y=35885
X2907 140 101 71 71 101 INV_X1 $T=65600 34600 1 0 $X=65485 $Y=33085
X2908 139 101 71 69 101 INV_X1 $T=67690 37400 1 0 $X=67575 $Y=35885
X2909 97 101 71 79 101 INV_X1 $T=68260 37400 1 0 $X=68145 $Y=35885
X3037 353 192 71 253 31 24 101 252 248 AOI222_X1 $T=21900 40200 0 180 $X=20265 $Y=38685
X3038 156 29 71 184 32 33 101 187 251 AOI222_X1 $T=20380 40200 0 0 $X=20265 $Y=40085
X3039 119 259 71 46 39 49 101 315 181 AOI222_X1 $T=34820 34600 0 0 $X=34705 $Y=34485
X3040 127 45 71 47 48 50 101 210 122 AOI222_X1 $T=35010 34600 1 0 $X=34895 $Y=33085
X3041 127 264 71 45 48 51 101 317 190 AOI222_X1 $T=36910 37400 1 0 $X=36795 $Y=35885
X3042 127 262 71 52 48 50 101 263 211 AOI222_X1 $T=38430 34600 1 0 $X=38315 $Y=33085
X3043 127 52 71 264 48 51 101 294 101 AOI222_X1 $T=40330 37400 0 0 $X=40215 $Y=37285
X3044 127 265 71 262 48 51 101 340 327 AOI222_X1 $T=40710 37400 1 0 $X=40595 $Y=35885
X3045 127 55 71 265 48 51 101 341 316 AOI222_X1 $T=42230 37400 1 0 $X=42115 $Y=35885
X3046 127 57 71 55 48 51 101 342 356 AOI222_X1 $T=45650 40200 0 180 $X=44015 $Y=38685
X3047 93 59 71 60 87 61 101 205 330 AOI222_X1 $T=47550 37400 1 0 $X=47435 $Y=35885
X3048 133 91 71 92 61 93 101 97 279 AOI222_X1 $T=62370 37400 0 0 $X=62255 $Y=37285
X3049 138 94 71 95 96 98 101 91 337 AOI222_X1 $T=64080 34600 0 0 $X=63965 $Y=34485
X3050 93 92 71 72 61 98 101 95 304 AOI222_X1 $T=67690 37400 0 180 $X=66055 $Y=35885
X3051 93 99 71 65 87 61 101 62 214 AOI222_X1 $T=67500 34600 0 0 $X=67385 $Y=34485
X3052 93 72 71 99 87 61 101 65 357 AOI222_X1 $T=67500 37400 0 0 $X=67385 $Y=37285
X3053 87 101 71 97 74 71 101 91 305 AOI222_X1 $T=67880 40200 0 0 $X=67765 $Y=40085
X3076 49 17 6 101 71 DLH_X1 $T=4230 37400 1 0 $X=4115 $Y=35885
X3077 49 21 7 101 71 DLH_X1 $T=7080 34600 0 0 $X=6965 $Y=34485
X3078 49 198 38 101 71 DLH_X1 $T=29500 40200 1 180 $X=27485 $Y=40085
X3079 49 200 39 101 71 DLH_X1 $T=29500 40200 0 0 $X=29385 $Y=40085
X3080 49 188 40 101 71 DLH_X1 $T=32160 37400 0 180 $X=30145 $Y=35885
X3081 49 201 259 101 71 DLH_X1 $T=32540 40200 1 0 $X=32425 $Y=38685
X3082 120 121 44 101 71 DLH_X1 $T=33870 37400 0 0 $X=33755 $Y=37285
X3083 50 202 264 101 71 DLH_X1 $T=39950 34600 1 0 $X=39835 $Y=33085
X3084 51 203 262 101 71 DLH_X1 $T=39950 34600 0 0 $X=39835 $Y=34485
X3085 128 263 267 101 71 DLH_X1 $T=42230 34600 1 0 $X=42115 $Y=33085
X3086 51 205 265 101 71 DLH_X1 $T=44130 40200 0 180 $X=42115 $Y=38685
X3087 128 317 56 101 71 DLH_X1 $T=42800 34600 0 0 $X=42685 $Y=34485
X3088 51 60 55 101 71 DLH_X1 $T=43750 37400 1 0 $X=43635 $Y=35885
X3089 128 341 58 101 71 DLH_X1 $T=44700 34600 0 0 $X=44585 $Y=34485
X3090 128 340 268 101 71 DLH_X1 $T=45650 37400 1 0 $X=45535 $Y=35885
X3091 128 294 269 101 71 DLH_X1 $T=45650 40200 1 0 $X=45535 $Y=38685
X3092 51 62 64 101 71 DLH_X1 $T=49070 40200 0 0 $X=48955 $Y=40085
X3093 51 59 57 101 71 DLH_X1 $T=49260 40200 1 0 $X=49145 $Y=38685
X3094 51 65 67 101 71 DLH_X1 $T=50970 40200 0 0 $X=50855 $Y=40085
X3095 128 342 66 101 71 DLH_X1 $T=53060 40200 0 180 $X=51045 $Y=38685
X3096 128 132 70 101 71 DLH_X1 $T=53060 40200 1 0 $X=52945 $Y=38685
X3097 51 139 75 101 71 DLH_X1 $T=57050 40200 1 180 $X=55035 $Y=40085
X3098 51 94 82 101 71 DLH_X1 $T=57050 40200 0 0 $X=56935 $Y=40085
X3099 38 39 43 42 101 71 118 OR4_X1 $T=33680 40200 1 180 $X=32425 $Y=40085
X3100 123 71 44 259 40 189 101 NOR4_X1 $T=36720 37400 1 180 $X=35655 $Y=37285
X3118 177 9 345 10 101 71 AOI21_X1 $T=8980 34600 1 0 $X=8865 $Y=33085
X3119 283 12 284 239 101 71 AOI21_X1 $T=11260 34600 0 0 $X=11145 $Y=34485
X3120 309 12 285 311 101 71 AOI21_X1 $T=11450 37400 1 0 $X=11335 $Y=35885
X3121 107 242 106 338 101 71 AOI21_X1 $T=13920 34600 1 180 $X=13045 $Y=34485
X3122 108 16 346 10 101 71 AOI21_X1 $T=15630 37400 0 180 $X=14755 $Y=35885
X3123 33 21 287 347 101 71 AOI21_X1 $T=17530 37400 1 0 $X=17415 $Y=35885
X3124 326 258 292 313 101 71 AOI21_X1 $T=28170 37400 1 180 $X=27295 $Y=37285
X3125 129 62 348 61 101 71 AOI21_X1 $T=48310 34600 1 0 $X=48195 $Y=33085
X3126 133 62 296 297 101 71 AOI21_X1 $T=51540 37400 0 180 $X=50665 $Y=35885
X3127 98 97 220 141 101 71 AOI21_X1 $T=65980 34600 1 0 $X=65865 $Y=33085
X3133 240 237 101 241 243 71 22 347 OAI221_X1 $T=12780 40200 1 0 $X=12665 $Y=38685
X3134 101 295 101 266 54 71 126 218 OAI221_X1 $T=41470 40200 0 0 $X=41355 $Y=40085
X3135 89 80 101 275 83 71 79 86 OAI221_X1 $T=60660 37400 1 180 $X=59405 $Y=37285
X3136 177 17 71 9 282 145 101 AOI22_X1 $T=7080 40200 0 180 $X=6015 $Y=38685
X3137 177 104 71 23 236 145 101 AOI22_X1 $T=8600 37400 0 0 $X=8485 $Y=37285
X3138 243 184 71 12 241 240 101 AOI22_X1 $T=11830 40200 1 0 $X=11715 $Y=38685
X3139 310 22 71 13 239 238 101 AOI22_X1 $T=13160 37400 0 180 $X=12095 $Y=35885
X3140 286 107 71 17 247 33 101 AOI22_X1 $T=13730 37400 0 0 $X=13615 $Y=37285
X3141 158 9 71 114 194 23 101 AOI22_X1 $T=20190 34600 0 180 $X=19125 $Y=33085
X3142 172 173 71 195 196 20 101 AOI22_X1 $T=24940 40200 1 180 $X=23875 $Y=40085
X3143 37 197 71 288 256 289 101 AOI22_X1 $T=25510 40200 0 180 $X=24445 $Y=38685
X3144 349 203 71 99 300 81 101 AOI22_X1 $T=58000 34600 1 180 $X=56935 $Y=34485
X3145 87 94 71 95 334 93 101 AOI22_X1 $T=57050 40200 1 0 $X=56935 $Y=38685
X3146 93 94 71 95 275 133 101 AOI22_X1 $T=58570 37400 0 0 $X=58455 $Y=37285
X3147 74 59 71 60 191 133 101 AOI22_X1 $T=58760 34600 1 0 $X=58645 $Y=33085
X3148 343 62 71 97 335 96 101 AOI22_X1 $T=60280 34600 1 180 $X=59215 $Y=34485
X3149 87 97 71 94 336 133 101 AOI22_X1 $T=60850 40200 1 180 $X=59785 $Y=40085
X3150 133 65 71 59 302 87 101 AOI22_X1 $T=61990 37400 0 180 $X=60925 $Y=35885
X3151 93 91 71 95 274 74 101 AOI22_X1 $T=61040 40200 1 0 $X=60925 $Y=38685
X3152 138 92 71 72 280 81 101 AOI22_X1 $T=62940 34600 0 180 $X=61875 $Y=33085
X3153 74 94 71 95 278 71 101 AOI22_X1 $T=61990 40200 1 0 $X=61875 $Y=38685
X3154 138 139 71 92 276 98 101 AOI22_X1 $T=62370 34600 0 0 $X=62255 $Y=34485
X3155 133 97 71 91 320 74 101 AOI22_X1 $T=64460 40200 1 180 $X=63395 $Y=40085
X3156 133 139 71 94 344 81 101 AOI22_X1 $T=65030 40200 0 0 $X=64915 $Y=40085
X3157 81 97 71 139 281 71 101 AOI22_X1 $T=65600 37400 0 0 $X=65485 $Y=37285
X3158 74 92 71 101 321 133 101 AOI22_X1 $T=69020 40200 0 180 $X=67955 $Y=38685
X3159 352 101 71 350 CLKBUF_X1 $T=1380 34600 0 0 $X=1265 $Y=34485
X3160 322 101 71 351 CLKBUF_X1 $T=2710 40200 0 0 $X=2595 $Y=40085
X3161 125 101 71 51 CLKBUF_X1 $T=39000 37400 0 180 $X=38315 $Y=35885
X3162 306 252 101 146 145 144 71 OAI22_X1 $T=2710 40200 1 180 $X=1645 $Y=40085
X3163 306 249 101 103 145 149 71 OAI22_X1 $T=5370 40200 0 0 $X=5255 $Y=40085
X3164 286 13 101 311 237 309 71 OAI22_X1 $T=12590 37400 1 180 $X=11525 $Y=37285
X3165 242 13 101 338 237 168 71 OAI22_X1 $T=12590 34600 1 0 $X=12475 $Y=33085
X3166 108 113 101 245 30 155 71 OAI22_X1 $T=16200 40200 0 0 $X=16085 $Y=40085
X3167 288 289 101 325 36 290 71 OAI22_X1 $T=23800 37400 1 0 $X=23685 $Y=35885
X3168 37 197 101 314 71 159 71 OAI22_X1 $T=27600 40200 1 180 $X=26535 $Y=40085
X3170 282 10 71 235 236 101 8 309 AOI221_X1 $T=9930 37400 1 0 $X=9815 $Y=35885
X3171 245 8 71 246 15 101 10 286 AOI221_X1 $T=13920 40200 1 0 $X=13805 $Y=38685
X3172 109 17 71 248 19 101 104 250 AOI221_X1 $T=16770 37400 0 0 $X=16655 $Y=37285
X3173 30 249 71 250 16 101 244 324 AOI221_X1 $T=17340 34600 0 0 $X=17225 $Y=34485
X3174 255 21 71 185 254 101 187 353 AOI221_X1 $T=21900 40200 1 0 $X=21785 $Y=38685
X3175 133 59 71 271 71 101 65 332 AOI221_X1 $T=53630 37400 1 0 $X=53515 $Y=35885
X3176 71 72 71 272 74 101 99 355 AOI221_X1 $T=55340 37400 0 0 $X=55225 $Y=37285
X3177 71 94 71 277 81 101 95 303 AOI221_X1 $T=62370 37400 1 0 $X=62255 $Y=35885
X3178 103 8 307 308 101 71 101 OAI21_X1 $T=8030 40200 0 0 $X=7915 $Y=40085
X3179 282 235 308 150 101 71 101 OAI21_X1 $T=8220 40200 1 0 $X=8105 $Y=38685
X3180 283 237 178 284 101 71 101 OAI21_X1 $T=10880 34600 1 0 $X=10765 $Y=33085
X3181 151 8 243 312 101 71 101 OAI21_X1 $T=12210 40200 0 0 $X=12095 $Y=40085
X3182 15 246 312 152 101 71 101 OAI21_X1 $T=14870 40200 0 0 $X=14755 $Y=40085
X3183 112 21 36 287 101 71 101 OAI21_X1 $T=20380 37400 0 180 $X=19505 $Y=35885
X3184 325 256 313 291 101 71 101 OAI21_X1 $T=24940 37400 0 0 $X=24825 $Y=37285
X3185 136 135 219 331 101 71 101 OAI21_X1 $T=56290 40200 0 180 $X=55415 $Y=38685
X3186 136 80 78 334 101 71 101 OAI21_X1 $T=56290 40200 1 0 $X=56175 $Y=38685
X3187 134 88 349 83 101 71 101 OAI21_X1 $T=57050 34600 1 0 $X=56935 $Y=33085
X3188 176 84 343 137 101 71 101 OAI21_X1 $T=59710 34600 1 0 $X=59595 $Y=33085
X3189 145 101 208 306 71 NAND2_X1 $T=3280 40200 1 0 $X=3165 $Y=38685
X3190 208 101 11 235 71 NAND2_X1 $T=8980 40200 1 0 $X=8865 $Y=38685
X3191 11 101 10 150 71 NAND2_X1 $T=9930 40200 1 0 $X=9815 $Y=38685
X3192 14 101 10 152 71 NAND2_X1 $T=15630 40200 0 180 $X=14945 $Y=38685
X3193 14 101 154 246 71 NAND2_X1 $T=15630 40200 0 0 $X=15515 $Y=40085
X3194 170 101 20 13 71 NAND2_X1 $T=17530 34600 1 0 $X=17415 $Y=33085
X3195 18 101 20 22 71 NAND2_X1 $T=19050 34600 1 180 $X=18365 $Y=34485
X3196 290 101 36 291 71 NAND2_X1 $T=24750 37400 1 0 $X=24635 $Y=35885
X3197 25 101 26 111 71 NAND2_X1 $T=36340 34600 0 0 $X=36225 $Y=34485
X3198 160 101 126 295 71 NAND2_X1 $T=38620 37400 0 0 $X=38505 $Y=37285
X3199 329 101 120 266 71 NAND2_X1 $T=43180 40200 1 180 $X=42495 $Y=40085
X3200 87 101 95 331 71 NAND2_X1 $T=54960 40200 1 0 $X=54845 $Y=38685
X3201 81 101 101 301 71 NAND2_X1 $T=56480 37400 0 0 $X=56365 $Y=37285
X3202 303 101 320 167 71 NAND2_X1 $T=62940 40200 0 0 $X=62825 $Y=40085
X3203 314 71 325 258 101 NOR2_X1 $T=27410 37400 1 180 $X=26725 $Y=37285
X3204 160 71 119 293 101 NOR2_X1 $T=31970 34600 0 0 $X=31855 $Y=34485
X3205 295 46 101 71 INV_X2 $T=40140 40200 1 0 $X=40025 $Y=38685
X3206 68 71 164 79 101 297 NOR3_X1 $T=52300 37400 0 180 $X=51425 $Y=35885
X3207 76 71 77 79 101 299 NOR3_X1 $T=56290 34600 1 0 $X=56175 $Y=33085
X3208 339 354 289 288 71 101 47 FA_X1 $T=24750 34600 0 0 $X=24635 $Y=34485
X3209 354 257 159 71 71 101 45 FA_X1 $T=25320 37400 1 0 $X=25205 $Y=35885
X3210 257 37 197 326 71 101 264 FA_X1 $T=25510 40200 1 0 $X=25395 $Y=38685
X3211 328 260 212 217 71 101 262 FA_X1 $T=37100 40200 1 0 $X=36985 $Y=38685
X3212 260 53 193 223 71 101 265 FA_X1 $T=38430 40200 0 0 $X=38315 $Y=40085
X3213 101 290 221 339 71 XNOR2_X1 $T=23610 34600 0 0 $X=23495 $Y=34485
X3214 101 215 261 328 71 XNOR2_X1 $T=34440 40200 1 0 $X=34325 $Y=38685
X3215 101 216 52 261 71 XNOR2_X1 $T=37480 37400 0 0 $X=37365 $Y=37285
X3218 112 17 285 71 247 101 101 OAI211_X1 $T=15630 37400 1 180 $X=14565 $Y=37285
X3219 32 22 171 71 251 288 101 OAI211_X1 $T=18290 40200 0 0 $X=18175 $Y=40085
X3220 140 63 330 71 296 318 101 OAI211_X1 $T=49070 34600 0 0 $X=48955 $Y=34485
X3221 83 69 336 71 274 165 101 OAI211_X1 $T=58950 40200 0 0 $X=58835 $Y=40085
X3222 83 85 302 71 276 273 101 OAI211_X1 $T=60090 37400 1 0 $X=59975 $Y=35885
X3223 89 69 278 71 279 166 101 OAI211_X1 $T=61040 37400 0 0 $X=60925 $Y=37285
X3224 111 109 101 24 25 26 71 252 27 OAI222_X1 $T=19430 37400 0 0 $X=19315 $Y=37285
X3225 111 158 101 16 25 26 71 244 28 OAI222_X1 $T=20190 34600 1 0 $X=20075 $Y=33085
X3226 111 19 101 30 25 26 71 249 34 OAI222_X1 $T=20380 34600 0 0 $X=20265 $Y=34485
X3227 111 255 101 31 25 26 71 253 290 OAI222_X1 $T=22280 37400 0 0 $X=22165 $Y=37285
X3228 111 254 101 35 25 26 71 29 289 OAI222_X1 $T=23040 40200 1 0 $X=22925 $Y=38685
X3229 137 69 101 88 83 89 71 90 277 OAI222_X1 $T=60470 34600 1 0 $X=60355 $Y=33085
X3230 236 10 235 101 345 283 71 AOI211_X1 $T=8980 34600 0 0 $X=8865 $Y=34485
X3231 10 244 169 101 235 168 71 AOI211_X1 $T=14490 34600 0 180 $X=13425 $Y=33085
X3232 245 10 246 101 346 310 71 AOI211_X1 $T=13920 37400 1 0 $X=13805 $Y=35885
X3233 10 158 153 101 246 242 71 AOI211_X1 $T=16200 34600 1 180 $X=15135 $Y=34485
X3234 33 23 157 101 184 179 71 AOI211_X1 $T=19430 34600 0 0 $X=19315 $Y=34485
X3235 74 65 318 101 270 298 71 AOI211_X1 $T=51540 34600 0 0 $X=51425 $Y=34485
X3236 98 72 73 101 299 333 71 AOI211_X1 $T=55340 34600 1 0 $X=55225 $Y=33085
X3239 183 157 18 101 71 NOR2_X2 $T=16580 34600 1 0 $X=16465 $Y=33085
X3240 61 74 213 101 71 NOR2_X2 $T=49070 34600 1 180 $X=48005 $Y=34485
X3241 131 101 175 280 298 267 71 NAND4_X1 $T=51160 34600 1 0 $X=51045 $Y=33085
X3242 333 101 300 206 332 269 71 NAND4_X1 $T=57050 37400 0 180 $X=55985 $Y=35885
X3243 335 101 301 319 355 268 71 NAND4_X1 $T=58000 37400 0 180 $X=56935 $Y=35885
X3244 281 101 321 337 357 207 71 NAND4_X1 $T=66550 37400 0 0 $X=66435 $Y=37285
X3246 84 164 69 101 90 163 68 271 71 OAI33_X1 $T=52110 34600 1 0 $X=51995 $Y=33085
X3247 84 77 80 101 69 163 134 270 71 OAI33_X1 $T=52490 34600 0 0 $X=52375 $Y=34485
X3248 80 134 164 101 77 68 135 272 71 OAI33_X1 $T=54770 37400 1 0 $X=54655 $Y=35885
X3249 116 101 224 174 71 199 NAND3_X1 $T=28930 34600 0 0 $X=28815 $Y=34485
X3250 305 101 344 304 71 222 NAND3_X1 $T=66740 40200 1 180 $X=65865 $Y=40085
X3252 293 120 101 71 BUF_X2 $T=32540 37400 0 0 $X=32425 $Y=37285
X3253 293 49 101 71 BUF_X2 $T=33110 37400 1 0 $X=32995 $Y=35885
X3256 115 101 71 2 CLKBUF_X3 $T=25130 40200 0 0 $X=25015 $Y=40085
X3257 41 101 71 4 CLKBUF_X3 $T=32160 37400 1 0 $X=32045 $Y=35885
.ENDS
***************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 10 A2 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 11 A3 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 8 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 A3 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS
** N=9 EP=5 IP=0 FDC=10
M0 6 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 9 A Z VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 8 A 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 7 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 7 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X2 VSS A B VDD ZN
** N=10 EP=5 IP=0 FDC=16
M0 6 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS 7 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 10 B VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=535 $Y=90 $D=1
M3 7 A 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=725 $Y=90 $D=1
M4 6 A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=1110 $Y=90 $D=1
M5 ZN A 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1300 $Y=90 $D=1
M6 6 B ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1490 $Y=90 $D=1
M7 ZN B 6 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1680 $Y=90 $D=1
M8 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M9 VDD 7 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M10 7 B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=535 $Y=680 $D=0
M11 VDD A 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=725 $Y=680 $D=0
M12 ZN A 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=1110 $Y=680 $D=0
M13 9 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1300 $Y=680 $D=0
M14 VDD B 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1490 $Y=680 $D=0
M15 8 B VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1680 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239
** N=397 EP=237 IP=4761 FDC=1816
M0 102 259 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=16385 $Y=29090 $D=1
M1 77 23 102 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16575 $Y=29090 $D=1
M2 102 23 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16765 $Y=29090 $D=1
M3 391 23 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=16940 $Y=26290 $D=1
M4 77 259 102 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16955 $Y=29090 $D=1
M5 27 106 391 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17130 $Y=26290 $D=1
M6 102 259 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17145 $Y=29090 $D=1
M7 392 106 27 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17320 $Y=26290 $D=1
M8 77 23 102 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17335 $Y=29090 $D=1
M9 77 23 392 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=17510 $Y=26290 $D=1
M10 102 23 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17525 $Y=29090 $D=1
M11 77 259 102 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=17715 $Y=29090 $D=1
M12 393 118 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=31165 $Y=31890 $D=1
M13 121 35 393 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31355 $Y=31890 $D=1
M14 394 35 121 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31545 $Y=31890 $D=1
M15 77 118 394 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31735 $Y=31890 $D=1
M16 395 31 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=31925 $Y=31890 $D=1
M17 121 267 395 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32115 $Y=31890 $D=1
M18 396 267 121 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=32305 $Y=31890 $D=1
M19 77 31 396 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=32495 $Y=31890 $D=1
M20 121 268 311 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=32870 $Y=31890 $D=1
M21 397 268 121 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33060 $Y=31890 $D=1
M22 77 29 397 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33250 $Y=31890 $D=1
M23 311 29 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=33440 $Y=31890 $D=1
M24 77 318 319 77 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=48645 $Y=31500 $D=1
M25 319 281 77 77 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=48835 $Y=31500 $D=1
M26 77 55 319 77 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=49025 $Y=31500 $D=1
M27 271 319 77 77 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=49215 $Y=31295 $D=1
M28 385 259 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=16385 $Y=29680 $D=0
M29 102 23 385 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16575 $Y=29680 $D=0
M30 386 23 102 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16765 $Y=29680 $D=0
M31 27 23 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=16940 $Y=26880 $D=0
M32 80 259 386 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16955 $Y=29680 $D=0
M33 80 106 27 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17130 $Y=26880 $D=0
M34 387 259 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17145 $Y=29680 $D=0
M35 27 106 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17320 $Y=26880 $D=0
M36 102 23 387 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17335 $Y=29680 $D=0
M37 80 23 27 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=17510 $Y=26880 $D=0
M38 388 23 102 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17525 $Y=29680 $D=0
M39 80 259 388 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=17715 $Y=29680 $D=0
M40 80 118 310 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=31165 $Y=32480 $D=0
M41 310 35 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31355 $Y=32480 $D=0
M42 80 35 310 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31545 $Y=32480 $D=0
M43 310 118 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31735 $Y=32480 $D=0
M44 312 31 310 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=31925 $Y=32480 $D=0
M45 310 267 312 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32115 $Y=32480 $D=0
M46 312 267 310 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=32305 $Y=32480 $D=0
M47 310 31 312 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=32495 $Y=32480 $D=0
M48 121 268 312 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=32870 $Y=32480 $D=0
M49 312 268 121 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33060 $Y=32480 $D=0
M50 121 29 312 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33250 $Y=32480 $D=0
M51 312 29 121 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=33440 $Y=32480 $D=0
M52 389 318 319 80 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=48645 $Y=30490 $D=0
M53 390 281 389 80 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=48835 $Y=30490 $D=0
M54 80 55 390 80 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=49025 $Y=30490 $D=0
M55 271 319 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=49215 $Y=30490 $D=0
X2331 379 6 77 80 10 77 DFF_X1 $T=1760 26200 0 0 $X=1645 $Y=26085
X2332 351 7 77 80 257 77 DFF_X1 $T=2330 29000 1 0 $X=2215 $Y=27485
X2333 352 6 77 80 256 77 DFF_X1 $T=2330 31800 1 0 $X=2215 $Y=30285
X2334 380 7 77 80 258 77 DFF_X1 $T=3090 26200 1 0 $X=2975 $Y=24685
X2335 303 6 77 80 34 77 DFF_X1 $T=26270 31800 1 0 $X=26155 $Y=30285
X2336 353 6 77 80 193 77 DFF_X1 $T=26270 31800 0 0 $X=26155 $Y=31685
X2337 340 6 77 80 32 77 DFF_X1 $T=28550 29000 1 0 $X=28435 $Y=27485
X2382 96 1 77 80 381 77 AND2_X1 $T=1000 26200 0 0 $X=885 $Y=26085
X2383 159 2 77 80 351 77 AND2_X1 $T=1190 29000 1 0 $X=1075 $Y=27485
X2384 96 3 77 80 339 77 AND2_X1 $T=1190 31800 1 0 $X=1075 $Y=30285
X2385 159 4 77 80 380 77 AND2_X1 $T=2330 26200 1 0 $X=2215 $Y=24685
X2386 159 5 77 80 160 77 AND2_X1 $T=2330 31800 0 0 $X=2215 $Y=31685
X2387 96 8 77 80 353 77 AND2_X1 $T=4990 31800 0 0 $X=4875 $Y=31685
X2388 96 9 77 80 340 77 AND2_X1 $T=7080 29000 1 0 $X=6965 $Y=27485
X2389 96 14 77 80 303 77 AND2_X1 $T=10120 31800 1 0 $X=10005 $Y=30285
X2390 273 50 77 80 316 77 AND2_X1 $T=43560 31800 1 0 $X=43445 $Y=30285
X2391 317 50 77 80 277 77 AND2_X1 $T=44320 31800 0 0 $X=44205 $Y=31685
X2392 317 275 77 80 136 77 AND2_X1 $T=45650 31800 0 0 $X=45535 $Y=31685
X2938 341 77 80 97 77 INV_X1 $T=8030 26200 1 180 $X=7535 $Y=26085
X2939 161 77 80 99 77 INV_X1 $T=10310 29000 0 0 $X=10195 $Y=28885
X2940 185 77 80 165 77 INV_X1 $T=16010 31800 0 180 $X=15515 $Y=30285
X2941 186 77 80 167 77 INV_X1 $T=16200 26200 1 0 $X=16085 $Y=24685
X2942 105 77 80 26 77 INV_X1 $T=17150 31800 0 180 $X=16655 $Y=30285
X2943 23 77 80 305 77 INV_X1 $T=17720 29000 1 0 $X=17605 $Y=27485
X2944 372 77 80 260 77 INV_X1 $T=20190 29000 0 180 $X=19695 $Y=27485
X2945 354 77 80 343 77 INV_X1 $T=20190 29000 1 0 $X=20075 $Y=27485
X2946 359 77 80 360 77 INV_X1 $T=25320 26200 1 0 $X=25205 $Y=24685
X2947 348 77 80 361 77 INV_X1 $T=27980 26200 1 180 $X=27485 $Y=26085
X2948 98 77 80 113 77 INV_X1 $T=32540 29000 1 180 $X=32045 $Y=28885
X2949 125 77 80 228 77 INV_X1 $T=34820 26200 1 0 $X=34705 $Y=24685
X2950 233 77 80 378 77 INV_X1 $T=36530 31800 1 0 $X=36415 $Y=30285
X2951 194 77 80 39 77 INV_X1 $T=38050 26200 0 0 $X=37935 $Y=26085
X2952 43 77 80 52 77 INV_X1 $T=40140 29000 0 0 $X=40025 $Y=28885
X2953 272 77 80 138 77 INV_X1 $T=41470 29000 0 180 $X=40975 $Y=27485
X2954 313 77 80 274 77 INV_X1 $T=41470 29000 1 0 $X=41355 $Y=27485
X2955 175 77 80 273 77 INV_X1 $T=42230 29000 1 0 $X=42115 $Y=27485
X2956 70 77 80 284 77 INV_X1 $T=50400 26200 0 180 $X=49905 $Y=24685
X2957 321 77 80 285 77 INV_X1 $T=50780 26200 1 180 $X=50285 $Y=26085
X2958 368 77 80 369 77 INV_X1 $T=57050 31800 1 0 $X=56935 $Y=30285
X2959 58 77 80 141 77 INV_X1 $T=61040 31800 0 0 $X=60925 $Y=31685
X2960 279 77 80 146 77 INV_X1 $T=62370 31800 0 0 $X=62255 $Y=31685
X2961 295 77 80 337 77 INV_X1 $T=63890 29000 0 0 $X=63775 $Y=28885
X2962 65 77 80 87 77 INV_X1 $T=65410 26200 1 180 $X=64915 $Y=26085
X2963 90 77 80 94 77 INV_X1 $T=68260 31800 0 180 $X=67765 $Y=30285
X2964 71 77 80 77 77 INV_X1 $T=68260 26200 0 0 $X=68145 $Y=26085
X3073 98 16 80 11 12 13 77 343 341 AOI222_X1 $T=9170 29000 1 0 $X=9055 $Y=27485
X3074 98 257 80 11 15 13 77 361 205 AOI222_X1 $T=9740 26200 0 0 $X=9625 $Y=26085
X3075 98 258 80 11 256 13 77 360 235 AOI222_X1 $T=11260 26200 1 0 $X=11145 $Y=24685
X3076 118 266 80 265 31 29 77 227 354 AOI222_X1 $T=29500 26200 1 180 $X=27865 $Y=26085
X3077 118 265 80 30 31 29 77 206 359 AOI222_X1 $T=29500 26200 1 0 $X=29385 $Y=24685
X3078 118 267 80 266 31 29 77 377 348 AOI222_X1 $T=29500 26200 0 0 $X=29385 $Y=26085
X3079 98 236 80 11 32 13 77 378 122 AOI222_X1 $T=32540 29000 0 0 $X=32425 $Y=28885
X3080 98 213 80 11 34 13 77 218 124 AOI222_X1 $T=33680 31800 0 0 $X=33565 $Y=31685
X3081 128 274 80 47 46 44 77 78 283 AOI222_X1 $T=45080 26200 1 180 $X=43445 $Y=26085
X3082 46 78 80 72 80 54 77 177 294 AOI222_X1 $T=58380 31800 1 0 $X=58265 $Y=30285
X3083 337 198 80 76 88 89 77 234 338 AOI222_X1 $T=65220 31800 1 0 $X=65105 $Y=30285
X3084 46 58 80 90 44 157 77 66 301 AOI222_X1 $T=69020 29000 0 180 $X=67385 $Y=27485
X3085 146 90 80 58 44 80 77 77 296 AOI222_X1 $T=69020 29000 1 180 $X=67385 $Y=28885
X3102 13 19 10 77 80 DLH_X1 $T=7650 29000 0 0 $X=7535 $Y=28885
X3103 13 21 256 77 80 DLH_X1 $T=9740 31800 1 180 $X=7725 $Y=31685
X3104 13 221 16 77 80 DLH_X1 $T=9740 31800 0 0 $X=9625 $Y=31685
X3105 13 216 17 77 80 DLH_X1 $T=11640 29000 1 0 $X=11525 $Y=27485
X3106 13 222 257 77 80 DLH_X1 $T=12400 29000 0 0 $X=12285 $Y=28885
X3107 13 103 258 77 80 DLH_X1 $T=14300 29000 0 0 $X=14185 $Y=28885
X3108 29 130 265 77 80 DLH_X1 $T=31020 26200 1 0 $X=30905 $Y=24685
X3109 29 133 266 77 80 DLH_X1 $T=33680 29000 0 180 $X=31665 $Y=27485
X3110 29 196 267 77 80 DLH_X1 $T=33680 29000 1 0 $X=33565 $Y=27485
X3111 29 47 35 77 80 DLH_X1 $T=38240 29000 1 180 $X=36225 $Y=28885
X3112 229 377 269 77 80 DLH_X1 $T=36720 26200 1 0 $X=36605 $Y=24685
X3113 29 78 36 77 80 DLH_X1 $T=37480 31800 0 0 $X=37365 $Y=31685
X3114 229 268 270 77 80 DLH_X1 $T=37860 29000 1 0 $X=37745 $Y=27485
X3115 29 194 37 77 80 DLH_X1 $T=38240 29000 0 0 $X=38125 $Y=28885
X3116 229 174 271 77 80 DLH_X1 $T=42610 31800 1 180 $X=40595 $Y=31685
X3117 15 80 12 256 10 347 77 NOR4_X1 $T=10690 29000 1 0 $X=10575 $Y=27485
X3118 257 80 16 258 17 100 77 NOR4_X1 $T=11260 26200 0 0 $X=11145 $Y=26085
X3119 177 80 49 278 133 382 77 NOR4_X1 $T=46220 29000 0 0 $X=46105 $Y=28885
X3120 60 80 62 282 323 365 77 NOR4_X1 $T=53060 26200 1 0 $X=52945 $Y=24685
X3121 152 80 67 79 150 336 77 NOR4_X1 $T=61990 26200 1 180 $X=60925 $Y=26085
X3139 102 21 342 215 77 80 AOI21_X1 $T=12400 31800 1 180 $X=11525 $Y=31685
X3140 110 261 372 345 77 80 AOI21_X1 $T=20570 29000 0 0 $X=20455 $Y=28885
X3141 314 40 363 133 77 80 AOI21_X1 $T=40330 29000 1 0 $X=40215 $Y=27485
X3142 284 49 45 315 77 80 AOI21_X1 $T=45080 26200 0 180 $X=44205 $Y=24685
X3143 53 214 280 39 77 80 AOI21_X1 $T=46220 26200 0 0 $X=46105 $Y=26085
X3144 74 278 318 51 77 80 AOI21_X1 $T=48500 31800 0 180 $X=47625 $Y=30285
X3145 65 77 142 324 77 80 AOI21_X1 $T=54390 31800 0 0 $X=54275 $Y=31685
X3146 144 53 326 51 77 80 AOI21_X1 $T=56480 26200 1 0 $X=56365 $Y=24685
X3147 145 292 368 141 77 80 AOI21_X1 $T=57620 29000 1 180 $X=56745 $Y=28885
X3148 80 82 374 336 77 80 AOI21_X1 $T=61990 29000 0 180 $X=61115 $Y=27485
X3153 109 169 77 27 28 80 115 114 OAI221_X1 $T=22280 31800 0 0 $X=22165 $Y=31685
X3154 199 91 77 286 287 80 152 269 OAI221_X1 $T=51920 26200 1 0 $X=51805 $Y=24685
X3155 74 77 77 299 87 80 64 298 OAI221_X1 $T=62370 26200 0 0 $X=62255 $Y=26085
X3156 153 91 77 300 279 80 67 181 OAI221_X1 $T=63510 31800 0 0 $X=63395 $Y=31685
X3157 295 51 77 301 87 80 93 375 OAI221_X1 $T=66360 29000 1 0 $X=66245 $Y=27485
X3158 166 163 80 19 304 102 77 AOI22_X1 $T=14870 31800 1 180 $X=13805 $Y=31685
X3159 217 162 80 18 164 119 77 AOI22_X1 $T=16200 26200 0 180 $X=15135 $Y=24685
X3160 105 169 80 224 306 108 77 AOI22_X1 $T=17910 31800 0 0 $X=17795 $Y=31685
X3161 77 225 80 356 262 112 77 AOI22_X1 $T=21900 31800 0 180 $X=20835 $Y=30285
X3162 46 82 80 72 299 157 77 AOI22_X1 $T=64460 26200 1 180 $X=63395 $Y=26085
X3163 63 77 80 66 302 44 77 AOI22_X1 $T=68450 31800 0 0 $X=68335 $Y=31685
X3164 381 77 80 379 CLKBUF_X1 $T=1380 26200 1 0 $X=1265 $Y=24685
X3165 339 77 80 352 CLKBUF_X1 $T=1380 29000 0 0 $X=1265 $Y=28885
X3166 264 77 80 98 CLKBUF_X1 $T=27220 29000 1 0 $X=27105 $Y=27485
X3167 33 77 80 29 CLKBUF_X1 $T=34440 26200 0 0 $X=34325 $Y=26085
X3168 356 112 77 344 308 114 80 OAI22_X1 $T=20950 29000 1 0 $X=20835 $Y=27485
X3169 77 225 77 355 358 173 80 OAI22_X1 $T=22280 31800 1 0 $X=22165 $Y=30285
X3170 53 200 77 293 126 74 80 OAI22_X1 $T=57240 26200 1 0 $X=57125 $Y=24685
X3177 364 40 80 280 54 77 43 383 AOI221_X1 $T=49260 26200 1 180 $X=48005 $Y=26085
X3178 80 49 80 289 63 77 177 366 AOI221_X1 $T=54200 29000 0 180 $X=52945 $Y=27485
X3179 86 57 80 85 84 77 77 287 AOI221_X1 $T=62940 26200 0 180 $X=61685 $Y=24685
X3180 297 68 80 298 77 77 148 371 AOI221_X1 $T=62180 29000 0 0 $X=62065 $Y=28885
X3181 63 183 80 375 54 77 77 300 AOI221_X1 $T=67880 31800 0 180 $X=66625 $Y=30285
X3182 26 20 223 184 77 80 77 OAI21_X1 $T=15630 31800 0 180 $X=14755 $Y=30285
X3183 111 21 358 342 77 80 77 OAI21_X1 $T=14870 31800 0 0 $X=14755 $Y=31685
X3184 169 24 211 104 77 80 77 OAI21_X1 $T=17910 31800 1 180 $X=17035 $Y=31685
X3185 305 260 187 185 77 80 77 OAI21_X1 $T=19050 29000 1 0 $X=18935 $Y=27485
X3186 111 26 308 172 77 80 77 OAI21_X1 $T=21140 31800 0 0 $X=21025 $Y=31685
X3187 344 262 345 307 77 80 77 OAI21_X1 $T=21330 29000 0 0 $X=21215 $Y=28885
X3188 363 39 207 362 77 80 77 OAI21_X1 $T=39190 26200 1 0 $X=39075 $Y=24685
X3189 382 276 132 82 77 80 77 OAI21_X1 $T=47360 29000 0 180 $X=46485 $Y=27485
X3190 290 57 364 135 77 80 77 OAI21_X1 $T=49640 29000 0 180 $X=48765 $Y=27485
X3191 75 77 332 53 77 80 77 OAI21_X1 $T=58000 29000 1 0 $X=57885 $Y=27485
X3192 67 90 231 64 77 80 77 OAI21_X1 $T=65980 26200 1 0 $X=65865 $Y=24685
X3193 107 77 25 161 80 NAND2_X1 $T=16390 29000 1 0 $X=16275 $Y=27485
X3194 259 77 305 111 80 NAND2_X1 $T=18480 29000 1 180 $X=17795 $Y=28885
X3195 171 77 170 20 80 NAND2_X1 $T=20190 26200 0 180 $X=19505 $Y=24685
X3196 114 77 308 307 80 NAND2_X1 $T=23230 29000 1 180 $X=22545 $Y=28885
X3197 39 77 176 313 80 NAND2_X1 $T=39190 26200 0 180 $X=38505 $Y=24685
X3198 384 77 195 362 80 NAND2_X1 $T=40520 26200 0 180 $X=39835 $Y=24685
X3199 39 77 41 272 80 NAND2_X1 $T=41280 26200 1 0 $X=41165 $Y=24685
X3200 317 77 273 127 80 NAND2_X1 $T=42230 29000 0 0 $X=42115 $Y=28885
X3201 78 77 52 42 80 NAND2_X1 $T=43560 26200 1 180 $X=42875 $Y=26085
X3202 316 77 314 288 80 NAND2_X1 $T=44510 29000 0 0 $X=44395 $Y=28885
X3203 274 77 316 129 80 NAND2_X1 $T=44890 29000 1 0 $X=44775 $Y=27485
X3204 316 77 317 152 80 NAND2_X1 $T=45080 31800 1 0 $X=44965 $Y=30285
X3205 277 77 48 219 80 NAND2_X1 $T=45080 31800 0 0 $X=44965 $Y=31685
X3206 131 77 130 53 80 NAND2_X1 $T=46410 26200 0 180 $X=45725 $Y=24685
X3207 275 77 47 135 80 NAND2_X1 $T=46410 31800 1 0 $X=46295 $Y=30285
X3208 275 77 277 180 80 NAND2_X1 $T=46410 31800 0 0 $X=46295 $Y=31685
X3209 277 77 134 81 80 NAND2_X1 $T=47740 31800 0 0 $X=47625 $Y=31685
X3210 316 77 138 290 80 NAND2_X1 $T=49640 29000 1 0 $X=49525 $Y=27485
X3211 333 77 322 281 80 NAND2_X1 $T=50400 31800 1 0 $X=50285 $Y=30285
X3212 177 77 51 92 80 NAND2_X1 $T=52300 31800 0 0 $X=52185 $Y=31685
X3213 68 77 66 144 80 NAND2_X1 $T=55910 26200 1 0 $X=55795 $Y=24685
X3214 201 77 148 147 80 NAND2_X1 $T=58950 26200 1 0 $X=58835 $Y=24685
X3215 44 77 177 370 80 NAND2_X1 $T=60280 29000 1 180 $X=59595 $Y=28885
X3216 203 77 76 209 80 NAND2_X1 $T=63510 26200 0 180 $X=62825 $Y=24685
X3217 68 77 148 295 80 NAND2_X1 $T=65220 29000 0 180 $X=64535 $Y=27485
X3218 77 77 77 335 80 NAND2_X1 $T=66360 26200 0 0 $X=66245 $Y=26085
X3219 165 80 106 166 77 NOR2_X1 $T=15630 31800 0 0 $X=15515 $Y=31685
X3220 185 80 306 259 77 NOR2_X1 $T=18480 31800 1 0 $X=18365 $Y=30285
X3221 355 80 344 261 77 NOR2_X1 $T=20380 31800 1 0 $X=20265 $Y=30285
X3222 188 80 357 226 77 NOR2_X1 $T=22850 26200 0 180 $X=22165 $Y=24685
X3223 31 80 123 33 77 NOR2_X1 $T=33870 26200 0 0 $X=33755 $Y=26085
X3224 47 80 196 314 77 NOR2_X1 $T=39760 29000 1 0 $X=39645 $Y=27485
X3225 272 80 47 317 77 NOR2_X1 $T=41280 29000 0 0 $X=41165 $Y=28885
X3226 78 80 43 50 77 NOR2_X1 $T=42990 31800 1 0 $X=42875 $Y=30285
X3227 197 80 130 275 77 NOR2_X1 $T=45270 26200 1 0 $X=45155 $Y=24685
X3228 288 80 51 276 77 NOR2_X1 $T=46030 29000 1 0 $X=45915 $Y=27485
X3229 292 80 46 65 77 NOR2_X1 $T=55530 29000 1 180 $X=54845 $Y=28885
X3230 180 80 83 77 77 NOR2_X1 $T=61420 31800 0 0 $X=61305 $Y=31685
X3231 92 80 152 89 77 NOR2_X1 $T=62370 31800 1 0 $X=62255 $Y=30285
X3232 152 80 51 88 77 NOR2_X1 $T=64270 26200 1 0 $X=64155 $Y=24685
X3233 272 80 175 52 77 315 NOR3_X1 $T=42230 26200 0 0 $X=42115 $Y=26085
X3234 288 80 83 94 77 349 NOR3_X1 $T=53060 31800 1 0 $X=52945 $Y=30285
X3235 64 80 83 290 77 291 NOR3_X1 $T=54200 29000 1 0 $X=54085 $Y=27485
X3236 129 80 143 93 77 324 NOR3_X1 $T=55910 31800 1 180 $X=55035 $Y=31685
X3237 94 80 129 156 77 327 NOR3_X1 $T=55910 31800 0 0 $X=55795 $Y=31685
X3238 325 80 291 326 77 331 NOR3_X1 $T=56290 29000 1 0 $X=56175 $Y=27485
X3239 70 80 147 79 77 330 NOR3_X1 $T=59710 26200 1 180 $X=58835 $Y=26085
X3240 373 263 112 356 80 77 30 FA_X1 $T=25320 29000 0 180 $X=22165 $Y=27485
X3241 263 346 173 358 80 77 265 FA_X1 $T=23230 29000 0 0 $X=23115 $Y=28885
X3242 346 77 225 110 80 77 266 FA_X1 $T=26270 31800 0 180 $X=23115 $Y=30285
X3243 77 162 185 18 80 XNOR2_X1 $T=13920 26200 0 180 $X=12665 $Y=24685
X3244 77 114 376 373 80 XNOR2_X1 $T=23420 26200 0 0 $X=23305 $Y=26085
X3245 77 308 123 376 80 XNOR2_X1 $T=25320 26200 0 180 $X=24065 $Y=24685
X3246 77 232 267 237 80 XNOR2_X1 $T=26270 31800 1 180 $X=25015 $Y=31685
X3247 111 19 304 80 101 356 77 OAI211_X1 $T=14870 31800 0 180 $X=13805 $Y=30285
X3248 335 81 202 80 294 328 77 OAI211_X1 $T=59710 31800 1 180 $X=58645 $Y=31685
X3249 149 126 370 80 374 350 77 OAI211_X1 $T=61230 29000 1 180 $X=60165 $Y=28885
X3250 149 61 371 80 296 151 77 OAI211_X1 $T=61230 29000 0 0 $X=61115 $Y=28885
X3251 279 64 338 80 154 182 77 OAI211_X1 $T=64650 31800 0 0 $X=64535 $Y=31685
X3252 153 94 204 80 302 155 77 OAI211_X1 $T=67500 31800 0 0 $X=67385 $Y=31685
X3253 131 39 77 52 53 279 80 56 282 OAI222_X1 $T=47740 26200 1 0 $X=47625 $Y=24685
X3254 156 93 77 67 92 91 80 51 297 OAI222_X1 $T=67500 29000 1 180 $X=65865 $Y=28885
X3255 139 43 349 77 367 322 80 AOI211_X1 $T=51350 31800 0 0 $X=51235 $Y=31685
X3256 146 71 328 77 327 329 80 AOI211_X1 $T=57620 31800 1 180 $X=56555 $Y=31685
X3257 63 72 330 77 293 220 80 AOI211_X1 $T=57050 29000 1 0 $X=56935 $Y=27485
X3258 332 78 350 77 334 333 80 AOI211_X1 $T=58760 29000 0 0 $X=58645 $Y=28885
X3265 158 77 148 316 138 137 80 NAND4_X1 $T=49450 29000 0 0 $X=49335 $Y=28885
X3266 329 77 369 73 331 178 80 NAND4_X1 $T=57430 31800 1 0 $X=57315 $Y=30285
X3267 148 77 64 94 77 210 80 NAND4_X1 $T=68070 26200 1 0 $X=67955 $Y=24685
X3269 189 190 191 77 117 116 309 264 80 OAI33_X1 $T=25700 26200 1 0 $X=25585 $Y=24685
X3270 52 313 200 77 272 42 126 384 80 OAI33_X1 $T=43560 26200 0 180 $X=42115 $Y=24685
X3271 59 290 156 77 92 129 61 367 80 OAI33_X1 $T=51730 31800 1 0 $X=51615 $Y=30285
X3272 141 290 92 77 156 288 61 289 80 OAI33_X1 $T=51920 29000 0 0 $X=51805 $Y=28885
X3273 77 92 288 77 75 83 61 321 80 OAI33_X1 $T=52490 26200 0 0 $X=52375 $Y=26085
X3274 94 143 75 77 70 83 59 323 80 OAI33_X1 $T=55150 26200 1 180 $X=53705 $Y=26085
X3275 143 288 91 77 67 69 70 325 80 OAI33_X1 $T=54960 29000 1 0 $X=54845 $Y=27485
X3276 290 143 67 77 93 69 288 238 80 OAI33_X1 $T=55720 31800 1 0 $X=55605 $Y=30285
X3277 64 143 70 77 295 179 59 334 80 OAI33_X1 $T=59710 26200 0 0 $X=59595 $Y=26085
X3278 20 77 168 167 80 25 NAND3_X1 $T=17340 26200 0 180 $X=16465 $Y=24685
X3279 24 77 171 170 80 107 NAND3_X1 $T=19620 26200 0 180 $X=18745 $Y=24685
X3280 306 77 165 305 80 109 NAND3_X1 $T=19810 31800 0 180 $X=18935 $Y=30285
X3281 347 77 192 212 80 309 NAND3_X1 $T=27600 26200 1 180 $X=26725 $Y=26085
X3282 314 77 273 194 80 153 NAND3_X1 $T=43750 29000 1 180 $X=42875 $Y=28885
X3283 273 77 314 177 80 214 NAND3_X1 $T=43370 29000 1 0 $X=43255 $Y=27485
X3284 315 77 48 176 80 279 NAND3_X1 $T=44320 26200 0 180 $X=43445 $Y=24685
X3285 58 77 277 134 80 278 NAND3_X1 $T=46980 31800 0 0 $X=46865 $Y=31685
X3286 136 77 78 52 80 292 NAND3_X1 $T=48690 29000 0 0 $X=48575 $Y=28885
X3287 198 77 284 58 80 320 NAND3_X1 $T=50020 26200 0 180 $X=49145 $Y=24685
X3288 140 77 365 366 80 270 NAND3_X1 $T=51730 26200 0 0 $X=51615 $Y=26085
X3289 239 77 76 56 80 208 NAND3_X1 $T=58190 26200 1 0 $X=58075 $Y=24685
X3291 38 77 80 230 CLKBUF_X3 $T=39380 31800 0 0 $X=39265 $Y=31685
X3292 283 285 320 383 77 80 286 AND4_X1 $T=49260 26200 0 0 $X=49145 $Y=26085
X3293 80 114 357 308 77 XOR2_X1 $T=21140 26200 1 0 $X=21025 $Y=24685
X3294 77 22 107 80 184 XNOR2_X2 $T=14870 26200 0 0 $X=14755 $Y=26085
X3295 77 25 22 80 104 XNOR2_X2 $T=20000 26200 0 0 $X=19885 $Y=26085
.ENDS
***************************************
.SUBCKT ICV_13
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6
** N=8 EP=6 IP=0 FDC=6
M0 7 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 93 94 95 96 97 98 99 100 101
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222
+ 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240 241 242
+ 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259
** N=465 EP=257 IP=5990 FDC=2084
M0 87 284 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=15815 $Y=22895 $D=1
M1 344 288 87 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16005 $Y=22895 $D=1
M2 87 288 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16195 $Y=22895 $D=1
M3 344 284 87 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16385 $Y=22895 $D=1
M4 87 284 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16575 $Y=22895 $D=1
M5 344 288 87 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16765 $Y=22895 $D=1
M6 87 288 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16955 $Y=22895 $D=1
M7 344 284 87 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17145 $Y=22895 $D=1
M8 53 343 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17335 $Y=22895 $D=1
M9 344 343 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17525 $Y=22895 $D=1
M10 53 343 344 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=17715 $Y=22895 $D=1
M11 344 343 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=17905 $Y=22895 $D=1
M12 94 350 352 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=22465 $Y=22895 $D=1
M13 352 288 94 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=22655 $Y=22895 $D=1
M14 94 288 352 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=22845 $Y=22895 $D=1
M15 352 350 94 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=23035 $Y=22895 $D=1
M16 53 351 352 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=23225 $Y=22895 $D=1
M17 352 351 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=23415 $Y=22895 $D=1
M18 103 353 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=28355 $Y=22895 $D=1
M19 53 353 103 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=28545 $Y=22895 $D=1
M20 463 21 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=28735 $Y=22895 $D=1
M21 353 27 463 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=28925 $Y=22895 $D=1
M22 109 302 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=37475 $Y=20690 $D=1
M23 53 302 109 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37665 $Y=20690 $D=1
M24 464 355 53 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37855 $Y=20690 $D=1
M25 109 29 464 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38045 $Y=20690 $D=1
M26 465 29 109 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38235 $Y=20690 $D=1
M27 53 355 465 53 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=38425 $Y=20690 $D=1
M28 457 284 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=15815 $Y=22090 $D=0
M29 87 288 457 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16005 $Y=22090 $D=0
M30 458 288 87 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16195 $Y=22090 $D=0
M31 80 284 458 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16385 $Y=22090 $D=0
M32 459 284 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16575 $Y=22090 $D=0
M33 87 288 459 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16765 $Y=22090 $D=0
M34 460 288 87 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16955 $Y=22090 $D=0
M35 80 284 460 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17145 $Y=22090 $D=0
M36 87 343 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17335 $Y=22090 $D=0
M37 80 343 87 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17525 $Y=22090 $D=0
M38 87 343 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=17715 $Y=22090 $D=0
M39 80 343 87 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=17905 $Y=22090 $D=0
M40 461 350 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=22465 $Y=22090 $D=0
M41 94 288 461 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=22655 $Y=22090 $D=0
M42 462 288 94 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=22845 $Y=22090 $D=0
M43 80 350 462 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=23035 $Y=22090 $D=0
M44 94 351 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=23225 $Y=22090 $D=0
M45 80 351 94 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=23415 $Y=22090 $D=0
M46 103 353 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=28355 $Y=22090 $D=0
M47 80 353 103 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=28545 $Y=22090 $D=0
M48 353 21 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=28735 $Y=22090 $D=0
M49 80 27 353 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=28925 $Y=22090 $D=0
M50 80 302 356 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=37475 $Y=21280 $D=0
M51 356 302 80 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37665 $Y=21280 $D=0
M52 109 355 356 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37855 $Y=21280 $D=0
M53 356 29 109 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38045 $Y=21280 $D=0
M54 109 29 356 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38235 $Y=21280 $D=0
M55 356 355 109 80 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=38425 $Y=21280 $D=0
X2876 402 3 53 80 152 53 DFF_X1 $T=1000 17800 0 0 $X=885 $Y=17685
X2877 449 3 53 80 228 53 DFF_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X2878 427 3 53 80 196 53 DFF_X1 $T=2330 20600 1 0 $X=2215 $Y=19085
X2879 452 3 53 80 151 53 DFF_X1 $T=5560 20600 1 180 $X=2215 $Y=20485
X2880 450 5 53 80 82 53 DFF_X1 $T=3090 17800 1 0 $X=2975 $Y=16285
X2881 426 5 53 80 7 53 DFF_X1 $T=4990 23400 1 0 $X=4875 $Y=21885
X2882 22 5 53 80 204 53 DFF_X1 $T=27220 20600 1 0 $X=27105 $Y=19085
X2883 249 5 53 80 173 53 DFF_X1 $T=34820 20600 1 0 $X=34705 $Y=19085
X2931 150 1 53 80 451 53 AND2_X1 $T=1190 15000 0 0 $X=1075 $Y=14885
X2932 195 2 53 80 450 53 AND2_X1 $T=2330 17800 1 0 $X=2215 $Y=16285
X2933 195 4 53 80 426 53 AND2_X1 $T=4230 23400 1 0 $X=4115 $Y=21885
X2934 81 273 53 80 452 53 AND2_X1 $T=6320 20600 1 180 $X=5445 $Y=20485
X2935 81 6 53 80 449 53 AND2_X1 $T=6700 23400 0 0 $X=6585 $Y=23285
X2936 81 274 53 80 402 53 AND2_X1 $T=7080 17800 0 0 $X=6965 $Y=17685
X2937 81 275 53 80 427 53 AND2_X1 $T=7080 20600 1 0 $X=6965 $Y=19085
X2938 10 9 53 80 276 53 AND2_X1 $T=10500 15000 1 180 $X=9625 $Y=14885
X2939 278 276 53 80 336 53 AND2_X1 $T=10310 20600 1 0 $X=10195 $Y=19085
X2940 81 26 53 80 171 53 AND2_X1 $T=35390 17800 1 180 $X=34515 $Y=17685
X2941 81 298 53 80 107 53 AND2_X1 $T=34820 15000 0 0 $X=34705 $Y=14885
X2942 81 299 53 80 243 53 AND2_X1 $T=35390 17800 0 0 $X=35275 $Y=17685
X2943 76 446 53 80 145 53 AND2_X1 $T=65410 23400 1 180 $X=64535 $Y=23285
X3608 153 53 80 273 53 INV_X1 $T=7460 23400 0 0 $X=7345 $Y=23285
X3609 13 53 80 217 53 INV_X1 $T=7840 15000 0 0 $X=7725 $Y=14885
X3610 439 53 80 274 53 INV_X1 $T=8600 20600 0 180 $X=8105 $Y=19085
X3611 428 53 80 333 53 INV_X1 $T=9360 17800 0 180 $X=8865 $Y=16285
X3612 250 53 80 275 53 INV_X1 $T=10310 23400 1 0 $X=10195 $Y=21885
X3613 9 53 80 337 53 INV_X1 $T=11070 15000 0 0 $X=10955 $Y=14885
X3614 342 53 80 279 53 INV_X1 $T=13540 20600 1 180 $X=13045 $Y=20485
X3615 156 53 80 239 53 INV_X1 $T=15440 23400 1 180 $X=14945 $Y=23285
X3616 444 53 80 283 53 INV_X1 $T=17340 20600 0 180 $X=16845 $Y=19085
X3617 86 53 80 407 53 INV_X1 $T=17150 15000 0 0 $X=17035 $Y=14885
X3618 163 53 80 286 53 INV_X1 $T=17530 15000 0 0 $X=17415 $Y=14885
X3619 165 53 80 345 53 INV_X1 $T=19810 20600 1 180 $X=19315 $Y=20485
X3620 90 53 80 411 53 INV_X1 $T=20570 15000 0 0 $X=20455 $Y=14885
X3621 409 53 80 231 53 INV_X1 $T=21330 23400 1 180 $X=20835 $Y=23285
X3622 290 53 80 410 53 INV_X1 $T=21140 15000 0 0 $X=21025 $Y=14885
X3623 93 53 80 347 53 INV_X1 $T=21900 23400 0 180 $X=21405 $Y=21885
X3624 349 53 80 348 53 INV_X1 $T=23040 17800 1 180 $X=22545 $Y=17685
X3625 287 53 80 16 53 INV_X1 $T=23990 17800 1 180 $X=23495 $Y=17685
X3626 289 53 80 412 53 INV_X1 $T=23990 23400 0 180 $X=23495 $Y=21885
X3627 95 53 80 97 53 INV_X1 $T=24940 20600 1 0 $X=24825 $Y=19085
X3628 291 53 80 440 53 INV_X1 $T=27030 15000 0 0 $X=26915 $Y=14885
X3629 415 53 80 23 53 INV_X1 $T=27980 20600 0 0 $X=27865 $Y=20485
X3630 24 53 80 292 53 INV_X1 $T=28170 23400 0 0 $X=28055 $Y=23285
X3631 89 53 80 96 53 INV_X1 $T=30450 20600 1 0 $X=30335 $Y=19085
X3632 105 53 80 298 53 INV_X1 $T=34250 20600 0 0 $X=34135 $Y=20485
X3633 106 53 80 299 53 INV_X1 $T=35390 23400 0 0 $X=35275 $Y=23285
X3634 172 53 80 32 53 INV_X1 $T=37670 23400 0 0 $X=37555 $Y=23285
X3635 174 53 80 176 53 INV_X1 $T=38050 23400 0 0 $X=37935 $Y=23285
X3636 30 53 80 31 53 INV_X1 $T=39570 17800 1 0 $X=39455 $Y=16285
X3637 359 53 80 37 53 INV_X1 $T=41470 23400 0 0 $X=41355 $Y=23285
X3638 175 53 80 36 53 INV_X1 $T=42230 20600 1 0 $X=42115 $Y=19085
X3639 305 53 80 111 53 INV_X1 $T=43180 20600 1 180 $X=42685 $Y=20485
X3640 420 53 80 221 53 INV_X1 $T=44700 17800 1 0 $X=44585 $Y=16285
X3641 69 53 80 42 53 INV_X1 $T=45080 17800 1 180 $X=44585 $Y=17685
X3642 366 53 80 308 53 INV_X1 $T=44890 23400 1 0 $X=44775 $Y=21885
X3643 44 53 80 67 53 INV_X1 $T=45840 17800 0 0 $X=45725 $Y=17685
X3644 116 53 80 117 53 INV_X1 $T=47930 20600 1 0 $X=47815 $Y=19085
X3645 33 53 80 311 53 INV_X1 $T=47930 20600 0 0 $X=47815 $Y=20485
X3646 123 53 80 66 53 INV_X1 $T=50780 20600 0 180 $X=50285 $Y=19085
X3647 212 53 80 118 53 INV_X1 $T=50780 20600 1 0 $X=50665 $Y=19085
X3648 49 53 80 127 53 INV_X1 $T=51730 17800 1 0 $X=51615 $Y=16285
X3649 436 53 80 377 53 INV_X1 $T=53250 20600 1 0 $X=53135 $Y=19085
X3650 320 53 80 316 53 INV_X1 $T=55150 17800 0 0 $X=55035 $Y=17685
X3651 129 53 80 178 53 INV_X1 $T=58190 15000 0 0 $X=58075 $Y=14885
X3652 382 53 80 323 53 INV_X1 $T=58380 20600 0 0 $X=58265 $Y=20485
X3653 136 53 80 190 53 INV_X1 $T=58570 15000 0 0 $X=58455 $Y=14885
X3654 60 53 80 149 53 INV_X1 $T=59520 15000 0 0 $X=59405 $Y=14885
X3655 326 53 80 70 53 INV_X1 $T=61040 17800 1 0 $X=60925 $Y=16285
X3656 192 53 80 223 53 INV_X1 $T=62180 15000 0 0 $X=62065 $Y=14885
X3657 396 53 80 324 53 INV_X1 $T=63320 17800 0 0 $X=63205 $Y=17685
X3658 325 53 80 328 53 INV_X1 $T=63700 20600 0 0 $X=63585 $Y=20485
X3659 45 53 80 125 53 INV_X1 $T=64650 17800 0 180 $X=64155 $Y=16285
X3660 77 53 80 236 53 INV_X1 $T=65980 15000 0 0 $X=65865 $Y=14885
X3661 147 53 80 48 53 INV_X1 $T=66360 17800 0 180 $X=65865 $Y=16285
X3662 424 53 80 51 53 INV_X1 $T=65980 23400 1 0 $X=65865 $Y=21885
X3663 148 53 80 246 53 INV_X1 $T=66740 15000 1 180 $X=66245 $Y=14885
X3664 126 53 80 248 53 INV_X1 $T=68070 17800 0 180 $X=67575 $Y=16285
X3665 143 53 80 53 53 INV_X1 $T=68070 17800 1 180 $X=67575 $Y=17685
X3666 400 53 80 331 53 INV_X1 $T=68260 15000 1 180 $X=67765 $Y=14885
X3667 58 53 80 79 53 INV_X1 $T=68070 17800 0 0 $X=67955 $Y=17685
X3668 53 53 80 57 53 INV_X1 $T=68450 20600 1 0 $X=68335 $Y=19085
X3790 229 7 80 8 11 12 53 447 439 AOI222_X1 $T=9360 23400 0 0 $X=9245 $Y=23285
X3810 12 230 13 53 80 DLH_X1 $T=13730 23400 0 180 $X=11715 $Y=21885
X3811 12 258 82 53 80 DLH_X1 $T=13160 23400 0 0 $X=13045 $Y=23285
X3812 12 158 15 53 80 DLH_X1 $T=13730 23400 1 0 $X=13615 $Y=21885
X3813 12 287 17 53 80 DLH_X1 $T=24180 17800 0 180 $X=22165 $Y=16285
X3814 12 289 18 53 80 DLH_X1 $T=23990 17800 0 0 $X=23875 $Y=17685
X3815 12 290 101 53 80 DLH_X1 $T=24180 17800 1 0 $X=24065 $Y=16285
X3816 12 409 19 53 80 DLH_X1 $T=24750 23400 0 0 $X=24635 $Y=23285
X3817 12 349 20 53 80 DLH_X1 $T=25320 20600 1 0 $X=25205 $Y=19085
X3818 206 416 24 53 80 DLH_X1 $T=28360 20600 0 0 $X=28245 $Y=20485
X3819 206 205 291 53 80 DLH_X1 $T=31970 17800 0 180 $X=29955 $Y=16285
X3820 109 295 296 53 80 DLH_X1 $T=30260 20600 0 0 $X=30145 $Y=20485
X3821 109 170 297 53 80 DLH_X1 $T=31400 23400 0 0 $X=31285 $Y=23285
X3822 109 294 25 53 80 DLH_X1 $T=31590 15000 0 0 $X=31475 $Y=14885
X3823 206 302 27 53 80 DLH_X1 $T=36340 23400 0 180 $X=34325 $Y=21885
X3824 109 433 300 53 80 DLH_X1 $T=35200 17800 1 0 $X=35085 $Y=16285
X3825 109 28 301 53 80 DLH_X1 $T=37670 23400 1 180 $X=35655 $Y=23285
X3826 163 80 157 289 290 430 53 NOR4_X1 $T=19050 17800 1 0 $X=18935 $Y=16285
X3827 19 80 18 20 101 413 53 NOR4_X1 $T=27790 17800 0 0 $X=27675 $Y=17685
X3828 303 80 417 108 416 355 53 NOR4_X1 $T=37480 17800 0 0 $X=37365 $Y=17685
X3829 57 80 58 436 63 379 53 NOR4_X1 $T=52300 20600 1 0 $X=52185 $Y=19085
X3830 64 80 65 62 382 187 53 NOR4_X1 $T=55340 23400 0 0 $X=55225 $Y=23285
X3856 334 279 253 403 53 80 AOI21_X1 $T=9550 20600 1 0 $X=9435 $Y=19085
X3857 277 10 334 337 53 80 AOI21_X1 $T=9740 17800 0 0 $X=9625 $Y=17685
X3858 405 278 428 404 53 80 AOI21_X1 $T=10880 17800 0 180 $X=10005 $Y=16285
X3859 84 14 339 337 53 80 AOI21_X1 $T=13730 15000 1 180 $X=12855 $Y=14885
X3860 103 292 447 354 53 80 AOI21_X1 $T=28550 23400 0 0 $X=28435 $Y=23285
X3861 21 295 354 27 53 80 AOI21_X1 $T=29120 23400 1 0 $X=29005 $Y=21885
X3862 174 32 360 207 53 80 AOI21_X1 $T=40710 17800 0 180 $X=39835 $Y=16285
X3863 454 305 361 445 53 80 AOI21_X1 $T=41850 20600 1 180 $X=40975 $Y=20485
X3864 306 37 307 363 53 80 AOI21_X1 $T=41660 23400 1 0 $X=41545 $Y=21885
X3865 221 42 421 222 53 80 AOI21_X1 $T=44700 15000 0 0 $X=44585 $Y=14885
X3866 235 44 369 174 53 80 AOI21_X1 $T=45080 17800 0 0 $X=44965 $Y=17685
X3867 122 52 120 396 53 80 AOI21_X1 $T=50400 15000 0 0 $X=50285 $Y=14885
X3868 113 37 124 245 53 80 AOI21_X1 $T=50970 17800 1 0 $X=50855 $Y=16285
X3869 251 50 441 396 53 80 AOI21_X1 $T=53060 15000 1 180 $X=52185 $Y=14885
X3870 378 319 213 45 53 80 AOI21_X1 $T=54010 20600 1 180 $X=53135 $Y=20485
X3871 379 61 319 383 53 80 AOI21_X1 $T=54390 20600 1 0 $X=54275 $Y=19085
X3872 381 227 386 147 53 80 AOI21_X1 $T=55720 15000 0 0 $X=55605 $Y=14885
X3873 386 68 385 123 53 80 AOI21_X1 $T=57430 15000 0 0 $X=57315 $Y=14885
X3874 137 50 442 78 53 80 AOI21_X1 $T=58950 23400 0 0 $X=58835 $Y=23285
X3875 146 72 224 225 53 80 AOI21_X1 $T=63510 15000 0 0 $X=63395 $Y=14885
X3876 397 79 443 140 53 80 AOI21_X1 $T=67690 20600 1 0 $X=67575 $Y=19085
X3877 59 79 401 53 53 80 AOI21_X1 $T=69020 23400 1 180 $X=68145 $Y=23285
X3880 38 112 53 307 40 80 67 366 OAI221_X1 $T=43750 23400 0 0 $X=43635 $Y=23285
X3881 369 46 53 41 309 80 436 114 OAI221_X1 $T=47170 15000 0 0 $X=47055 $Y=14885
X3882 148 194 53 331 77 80 252 247 OAI221_X1 $T=66740 15000 0 0 $X=66625 $Y=14885
X3883 281 278 80 282 280 338 53 AOI22_X1 $T=13730 20600 1 0 $X=13615 $Y=19085
X3884 84 14 80 159 342 157 53 AOI22_X1 $T=14680 15000 0 0 $X=14565 $Y=14885
X3885 339 341 80 159 240 157 53 AOI22_X1 $T=15060 17800 1 0 $X=14945 $Y=16285
X3886 429 444 80 86 404 286 53 AOI22_X1 $T=16010 17800 1 0 $X=15895 $Y=16285
X3887 286 86 80 407 444 163 53 AOI22_X1 $T=16960 17800 1 0 $X=16845 $Y=16285
X3888 96 407 80 286 226 89 53 AOI22_X1 $T=18480 15000 0 0 $X=18365 $Y=14885
X3889 89 164 80 241 415 96 53 AOI22_X1 $T=19810 23400 1 180 $X=18745 $Y=23285
X3890 412 93 80 347 165 289 53 AOI22_X1 $T=20760 20600 1 180 $X=19695 $Y=20485
X3891 410 90 80 411 285 290 53 AOI22_X1 $T=20950 17800 1 0 $X=20835 $Y=16285
X3892 453 285 80 411 431 290 53 AOI22_X1 $T=21900 17800 1 180 $X=20835 $Y=17685
X3893 348 287 80 16 288 349 53 AOI22_X1 $T=22850 20600 1 0 $X=22735 $Y=19085
X3894 89 412 80 347 199 96 53 AOI22_X1 $T=23420 20600 0 0 $X=23305 $Y=20485
X3895 103 23 80 433 432 206 53 AOI22_X1 $T=32920 17800 0 180 $X=31855 $Y=16285
X3896 365 235 80 44 418 434 53 AOI22_X1 $T=43180 20600 1 0 $X=43065 $Y=19085
X3897 455 147 80 37 422 184 53 AOI22_X1 $T=48880 23400 1 180 $X=47815 $Y=23285
X3898 423 108 80 44 121 310 53 AOI22_X1 $T=49640 23400 0 0 $X=49525 $Y=23285
X3899 135 42 80 191 392 323 53 AOI22_X1 $T=58760 23400 1 0 $X=58645 $Y=21885
X3900 443 53 80 48 332 425 53 AOI22_X1 $T=67120 20600 0 0 $X=67005 $Y=20485
X3901 451 53 80 238 CLKBUF_X1 $T=2330 15000 0 0 $X=2215 $Y=14885
X3902 279 337 53 338 155 83 80 OAI22_X1 $T=12970 15000 1 180 $X=11905 $Y=14885
X3903 283 431 53 282 86 286 80 OAI22_X1 $T=16200 17800 0 0 $X=16085 $Y=17685
X3904 88 345 53 284 347 289 80 OAI22_X1 $T=18670 23400 1 0 $X=18555 $Y=21885
X3905 345 166 53 350 93 412 80 OAI22_X1 $T=19620 23400 1 0 $X=19505 $Y=21885
X3906 96 410 53 168 411 89 80 OAI22_X1 $T=21520 15000 0 0 $X=21405 $Y=14885
X3907 96 348 53 169 16 89 80 OAI22_X1 $T=24750 15000 1 180 $X=23685 $Y=14885
X3908 98 201 53 99 414 80 80 OAI22_X1 $T=25510 20600 0 0 $X=25395 $Y=20485
X3909 369 46 53 419 174 43 80 OAI22_X1 $T=46220 17800 0 180 $X=45155 $Y=16285
X3910 34 36 53 310 53 45 80 OAI22_X1 $T=48310 23400 1 0 $X=48195 $Y=21885
X3911 143 216 53 400 215 126 80 OAI22_X1 $T=69020 17800 0 180 $X=67955 $Y=16285
X3918 279 154 80 280 281 53 341 254 AOI221_X1 $T=12590 20600 1 0 $X=12475 $Y=19085
X3919 440 202 80 21 291 53 234 293 AOI221_X1 $T=27410 15000 0 0 $X=27295 $Y=14885
X3920 206 294 80 293 103 53 291 203 AOI221_X1 $T=29690 15000 1 180 $X=28435 $Y=14885
X3921 304 177 80 34 362 53 176 445 AOI221_X1 $T=40520 23400 1 0 $X=40405 $Y=21885
X3922 358 360 80 35 437 53 110 456 AOI221_X1 $T=40710 17800 1 0 $X=40595 $Y=16285
X3923 312 175 80 313 314 53 125 371 AOI221_X1 $T=49830 23400 1 0 $X=49715 $Y=21885
X3924 441 52 80 315 55 53 61 309 AOI221_X1 $T=52300 15000 1 180 $X=51045 $Y=14885
X3925 123 67 80 69 316 53 384 321 AOI221_X1 $T=57430 17800 1 180 $X=56175 $Y=17685
X3926 333 276 335 277 53 80 53 OAI21_X1 $T=8980 17800 0 0 $X=8865 $Y=17685
X3927 334 279 403 335 53 80 53 OAI21_X1 $T=9930 20600 0 0 $X=9815 $Y=20485
X3928 349 16 408 343 53 80 53 OAI21_X1 $T=18290 20600 0 180 $X=17415 $Y=19085
X3929 408 285 255 346 53 80 53 OAI21_X1 $T=18480 17800 0 0 $X=18365 $Y=17685
X3930 290 411 429 346 53 80 53 OAI21_X1 $T=20000 17800 1 180 $X=19125 $Y=17685
X3931 348 287 453 351 53 80 53 OAI21_X1 $T=22850 20600 0 180 $X=21975 $Y=19085
X3932 21 23 219 432 53 80 53 OAI21_X1 $T=28740 17800 1 0 $X=28625 $Y=16285
X3933 43 30 358 32 53 80 53 OAI21_X1 $T=38240 17800 1 0 $X=38125 $Y=16285
X3934 360 31 363 357 53 80 53 OAI21_X1 $T=40330 17800 1 180 $X=39455 $Y=17685
X3935 418 33 296 361 53 80 53 OAI21_X1 $T=40330 20600 0 0 $X=40215 $Y=20485
X3936 207 36 454 32 53 80 53 OAI21_X1 $T=41090 20600 1 0 $X=40975 $Y=19085
X3937 42 39 434 41 53 80 53 OAI21_X1 $T=44890 20600 0 180 $X=44015 $Y=19085
X3938 113 41 435 32 53 80 53 OAI21_X1 $T=45080 20600 1 180 $X=44205 $Y=20485
X3939 34 47 312 115 53 80 53 OAI21_X1 $T=48310 23400 0 180 $X=47435 $Y=21885
X3940 46 48 315 66 53 80 53 OAI21_X1 $T=48880 17800 1 0 $X=48765 $Y=16285
X3941 49 48 423 116 53 80 53 OAI21_X1 $T=49640 23400 1 180 $X=48765 $Y=23285
X3942 143 56 455 374 53 80 53 OAI21_X1 $T=51730 23400 0 0 $X=51615 $Y=23285
X3943 79 147 384 53 53 80 53 OAI21_X1 $T=55530 17800 0 0 $X=55415 $Y=17685
X3944 322 321 365 387 53 80 53 OAI21_X1 $T=58760 17800 1 180 $X=57885 $Y=17685
X3945 392 48 394 388 53 80 53 OAI21_X1 $T=61040 20600 0 180 $X=60165 $Y=19085
X3946 134 48 142 144 53 80 53 OAI21_X1 $T=62370 23400 0 0 $X=62255 $Y=23285
X3947 401 78 399 398 53 80 53 OAI21_X1 $T=68260 23400 1 180 $X=67385 $Y=23285
X3948 9 53 154 405 80 NAND2_X1 $T=10500 15000 0 0 $X=10385 $Y=14885
X3949 404 53 336 277 80 NAND2_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X3950 83 53 155 278 80 NAND2_X1 $T=12020 17800 1 0 $X=11905 $Y=16285
X3951 282 53 278 340 80 NAND2_X1 $T=13540 17800 1 180 $X=12855 $Y=17685
X3952 340 53 10 341 80 NAND2_X1 $T=13540 17800 0 0 $X=13425 $Y=17685
X3953 84 53 159 291 80 NAND2_X1 $T=15630 15000 0 0 $X=15515 $Y=14885
X3954 160 53 162 241 80 NAND2_X1 $T=16390 23400 0 0 $X=16275 $Y=23285
X3955 284 53 288 343 80 NAND2_X1 $T=18670 23400 0 180 $X=17985 $Y=21885
X3956 408 53 285 346 80 NAND2_X1 $T=18290 20600 1 0 $X=18175 $Y=19085
X3957 350 53 288 351 80 NAND2_X1 $T=23610 23400 1 180 $X=22925 $Y=23285
X3958 108 53 176 304 80 NAND2_X1 $T=39000 23400 1 180 $X=38315 $Y=23285
X3959 115 53 32 359 80 NAND2_X1 $T=39000 23400 0 0 $X=38885 $Y=23285
X3960 115 53 31 305 80 NAND2_X1 $T=39760 20600 0 0 $X=39645 $Y=20485
X3961 39 53 36 362 80 NAND2_X1 $T=40900 23400 0 0 $X=40785 $Y=23285
X3962 111 53 176 364 80 NAND2_X1 $T=42800 20600 1 180 $X=42115 $Y=20485
X3963 36 53 31 113 80 NAND2_X1 $T=42990 17800 1 180 $X=42305 $Y=17685
X3964 111 53 32 34 80 NAND2_X1 $T=43750 20600 0 0 $X=43635 $Y=20485
X3965 37 53 30 116 80 NAND2_X1 $T=48120 17800 1 180 $X=47435 $Y=17685
X3966 311 53 47 49 80 NAND2_X1 $T=49640 20600 1 180 $X=48955 $Y=20485
X3967 311 53 41 56 80 NAND2_X1 $T=49260 23400 1 0 $X=49145 $Y=21885
X3968 119 53 138 436 80 NAND2_X1 $T=50400 20600 0 180 $X=49715 $Y=19085
X3969 119 53 135 126 80 NAND2_X1 $T=51730 20600 1 0 $X=51615 $Y=19085
X3970 376 53 50 122 80 NAND2_X1 $T=53630 15000 1 180 $X=52945 $Y=14885
X3971 316 53 66 317 80 NAND2_X1 $T=53440 17800 0 0 $X=53325 $Y=17685
X3972 380 53 377 186 80 NAND2_X1 $T=54960 23400 0 180 $X=54275 $Y=21885
X3973 324 53 50 62 80 NAND2_X1 $T=55720 20600 0 180 $X=55035 $Y=19085
X3974 119 53 66 382 80 NAND2_X1 $T=55720 20600 0 0 $X=55605 $Y=20485
X3975 54 53 42 134 80 NAND2_X1 $T=56860 23400 1 0 $X=56745 $Y=21885
X3976 78 53 57 129 80 NAND2_X1 $T=57810 23400 1 180 $X=57125 $Y=23285
X3977 54 53 119 326 80 NAND2_X1 $T=57430 17800 0 0 $X=57315 $Y=17685
X3978 377 53 123 148 80 NAND2_X1 $T=58760 20600 0 180 $X=58075 $Y=19085
X3979 190 53 70 60 80 NAND2_X1 $T=58950 15000 0 0 $X=58835 $Y=14885
X3980 138 53 67 320 80 NAND2_X1 $T=58950 17800 1 0 $X=58835 $Y=16285
X3981 380 53 70 214 80 NAND2_X1 $T=61040 15000 0 0 $X=60925 $Y=14885
X3982 70 53 147 77 80 NAND2_X1 $T=61420 17800 1 0 $X=61305 $Y=16285
X3983 70 53 50 325 80 NAND2_X1 $T=61990 23400 0 180 $X=61305 $Y=21885
X3984 125 53 70 192 80 NAND2_X1 $T=62180 15000 1 180 $X=61495 $Y=14885
X3985 71 53 48 136 80 NAND2_X1 $T=62370 17800 1 0 $X=62255 $Y=16285
X3986 53 53 53 327 80 NAND2_X1 $T=62940 17800 1 180 $X=62255 $Y=17685
X3987 324 53 191 68 80 NAND2_X1 $T=64270 23400 0 180 $X=63585 $Y=21885
X3988 53 53 48 396 80 NAND2_X1 $T=65410 17800 1 0 $X=65295 $Y=16285
X3989 76 53 57 74 80 NAND2_X1 $T=65980 20600 1 0 $X=65865 $Y=19085
X3990 57 53 79 424 80 NAND2_X1 $T=66550 20600 0 0 $X=66435 $Y=20485
X3991 279 80 337 281 53 NOR2_X1 $T=12970 17800 1 180 $X=12285 $Y=17685
X3992 160 80 158 197 53 NOR2_X1 $T=16390 23400 1 180 $X=15705 $Y=23285
X3993 91 80 409 167 53 NOR2_X1 $T=21330 23400 0 0 $X=21215 $Y=23285
X3994 364 80 39 110 53 NOR2_X1 $T=42800 17800 0 180 $X=42115 $Y=16285
X3995 123 80 135 54 53 NOR2_X1 $T=51160 20600 1 0 $X=51045 $Y=19085
X3996 62 80 64 380 53 NOR2_X1 $T=54960 23400 1 0 $X=54845 $Y=21885
X3997 21 104 53 80 INV_X2 $T=29500 17800 1 0 $X=29385 $Y=16285
X3998 69 80 108 181 53 220 NOR3_X1 $T=43750 17800 1 180 $X=42875 $Y=17685
X3999 39 80 174 30 53 375 NOR3_X1 $T=46790 17800 0 0 $X=46675 $Y=17685
X4000 126 80 49 53 53 313 NOR3_X1 $T=51730 23400 0 180 $X=50855 $Y=21885
X4001 62 80 129 59 53 318 NOR3_X1 $T=53060 17800 1 0 $X=52945 $Y=16285
X4002 130 80 58 71 53 381 NOR3_X1 $T=54770 17800 1 0 $X=54655 $Y=16285
X4003 325 80 58 71 53 29 NOR3_X1 $T=63130 20600 1 180 $X=62255 $Y=20485
X4004 53 283 218 429 80 XNOR2_X1 $T=15060 20600 1 0 $X=14945 $Y=19085
X4005 53 431 256 444 80 XNOR2_X1 $T=21140 20600 0 180 $X=19885 $Y=19085
X4006 53 285 232 453 80 XNOR2_X1 $T=20760 20600 0 0 $X=20645 $Y=20485
X4007 53 259 233 27 80 XNOR2_X1 $T=24750 23400 1 180 $X=23495 $Y=23285
X4009 367 45 370 80 308 297 53 OAI211_X1 $T=46030 20600 1 180 $X=44965 $Y=20485
X4010 385 320 41 80 143 437 53 OAI211_X1 $T=56480 17800 0 180 $X=55415 $Y=16285
X4011 332 325 389 80 390 314 53 OAI211_X1 $T=61420 23400 0 180 $X=60355 $Y=21885
X4012 147 42 438 53 135 322 80 AOI211_X1 $T=58000 17800 1 0 $X=57885 $Y=16285
X4013 327 50 123 53 69 438 80 AOI211_X1 $T=61040 17800 1 180 $X=59975 $Y=17685
X4014 391 50 326 53 327 393 80 AOI211_X1 $T=61040 17800 0 0 $X=60925 $Y=17685
X4015 395 328 394 53 393 367 80 AOI211_X1 $T=62940 20600 0 180 $X=61875 $Y=19085
X4016 329 74 396 53 75 448 80 AOI211_X1 $T=65220 17800 0 0 $X=65105 $Y=17685
X4017 237 57 75 53 58 425 80 AOI211_X1 $T=69020 20600 1 180 $X=67955 $Y=20485
X4021 302 115 416 53 80 NOR2_X2 $T=37290 23400 0 180 $X=36225 $Y=21885
X4022 342 53 336 406 161 85 80 NAND4_X1 $T=15820 20600 0 0 $X=15705 $Y=20485
X4023 430 53 348 83 198 91 80 NAND4_X1 $T=20000 17800 1 0 $X=19885 $Y=16285
X4024 200 53 80 413 100 414 80 NAND4_X1 $T=25320 23400 1 0 $X=25205 $Y=21885
X4025 19 53 18 20 101 242 80 NAND4_X1 $T=27790 17800 1 180 $X=26725 $Y=17685
X4026 177 53 32 66 42 211 80 NAND4_X1 $T=46220 17800 1 0 $X=46105 $Y=16285
X4027 422 53 368 183 371 301 80 NAND4_X1 $T=47930 23400 1 180 $X=46865 $Y=23285
X4028 375 53 48 75 140 303 80 NAND4_X1 $T=52680 17800 1 180 $X=51615 $Y=17685
X4029 70 53 324 127 73 133 80 NAND4_X1 $T=56290 20600 0 0 $X=56175 $Y=20485
X4030 188 53 380 54 42 189 80 NAND4_X1 $T=56290 23400 0 0 $X=56175 $Y=23285
X4034 304 43 30 53 175 47 176 306 80 OAI33_X1 $T=39190 23400 1 0 $X=39075 $Y=21885
X4035 209 364 47 53 138 180 421 210 80 OAI33_X1 $T=42230 15000 0 0 $X=42115 $Y=14885
X4036 362 359 138 53 66 112 34 179 80 OAI33_X1 $T=42420 23400 0 0 $X=42305 $Y=23285
X4037 42 33 39 53 53 45 135 372 80 OAI33_X1 $T=48500 20600 1 0 $X=48385 $Y=19085
X4038 128 420 69 53 317 373 303 185 80 OAI33_X1 $T=48690 17800 0 0 $X=48575 $Y=17685
X4039 63 62 374 53 49 60 75 131 80 OAI33_X1 $T=55340 23400 1 180 $X=53895 $Y=23285
X4040 140 134 136 53 317 68 75 383 80 OAI33_X1 $T=58190 20600 0 180 $X=56745 $Y=19085
X4041 141 129 391 53 140 382 68 257 80 OAI33_X1 $T=60660 23400 0 0 $X=60545 $Y=23285
X4042 53 320 123 53 63 424 325 446 80 OAI33_X1 $T=62370 23400 1 0 $X=62255 $Y=21885
X4043 78 79 147 53 76 65 391 330 80 OAI33_X1 $T=66740 23400 1 180 $X=65295 $Y=23285
X4044 358 53 115 175 80 357 NAND3_X1 $T=38810 20600 0 180 $X=37935 $Y=19085
X4045 419 53 36 31 80 208 NAND3_X1 $T=41850 15000 1 180 $X=40975 $Y=14885
X4046 178 53 177 32 80 417 NAND3_X1 $T=42420 17800 1 180 $X=41545 $Y=17685
X4047 43 53 32 182 80 420 NAND3_X1 $T=44700 17800 0 180 $X=43825 $Y=16285
X4048 435 53 115 174 80 368 NAND3_X1 $T=45270 23400 1 0 $X=45155 $Y=21885
X4049 372 53 123 67 80 370 NAND3_X1 $T=47930 20600 1 180 $X=47055 $Y=20485
X4050 222 53 51 50 80 373 NAND3_X1 $T=50400 17800 0 180 $X=49525 $Y=16285
X4051 318 53 375 316 80 128 NAND3_X1 $T=53440 17800 1 180 $X=52565 $Y=17685
X4052 57 53 59 79 80 376 NAND3_X1 $T=54390 15000 1 180 $X=53515 $Y=14885
X4053 130 53 29 188 80 378 NAND3_X1 $T=55720 20600 1 180 $X=54845 $Y=20485
X4054 79 53 61 323 80 139 NAND3_X1 $T=58760 20600 0 0 $X=58645 $Y=20485
X4055 377 53 190 58 80 388 NAND3_X1 $T=59520 20600 1 0 $X=59405 $Y=19085
X4056 323 53 190 53 80 389 NAND3_X1 $T=59520 20600 0 0 $X=59405 $Y=20485
X4057 442 53 377 324 80 390 NAND3_X1 $T=59710 23400 1 0 $X=59595 $Y=21885
X4058 178 53 73 48 80 397 NAND3_X1 $T=64460 17800 1 180 $X=63585 $Y=17685
X4059 140 53 51 73 80 329 NAND3_X1 $T=65220 17800 1 180 $X=64345 $Y=17685
X4060 399 53 324 328 80 387 NAND3_X1 $T=65220 20600 0 180 $X=64345 $Y=19085
X4061 324 53 59 79 80 391 NAND3_X1 $T=65220 23400 1 0 $X=65105 $Y=21885
X4062 193 53 51 132 80 398 NAND3_X1 $T=66740 23400 0 0 $X=66625 $Y=23285
X4064 285 288 444 165 53 80 406 AND4_X1 $T=17910 20600 1 180 $X=16655 $Y=20485
X4065 80 244 300 456 53 XOR2_X1 $T=38240 17800 0 180 $X=36985 $Y=16285
X4087 64 317 53 80 374 53 OR2_X1 $T=53440 23400 0 180 $X=52565 $Y=21885
X4088 448 330 53 80 395 53 OR2_X1 $T=65980 20600 0 180 $X=65105 $Y=19085
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7
** N=13 EP=7 IP=0 FDC=16
M0 12 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 12 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 9 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 9 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 13 A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 10 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 8 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 9 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 9 A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 10 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 10 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209
** N=387 EP=208 IP=4537 FDC=1902
M0 386 49 303 50 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=55865 $Y=6690 $D=1
M1 387 44 386 50 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=56055 $Y=6690 $D=1
M2 50 98 387 50 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=56245 $Y=6690 $D=1
M3 304 303 50 50 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=56435 $Y=6690 $D=1
M4 39 49 303 39 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=55865 $Y=7595 $D=0
M5 303 44 39 39 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=56055 $Y=7595 $D=0
M6 39 98 303 39 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=56245 $Y=7595 $D=0
M7 304 303 39 39 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=56435 $Y=7280 $D=0
X2145 340 4 50 39 115 50 DFF_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X2146 374 5 50 39 226 50 DFF_X1 $T=1760 9400 1 0 $X=1645 $Y=7885
X2147 375 5 50 39 223 50 DFF_X1 $T=2330 6600 0 0 $X=2215 $Y=6485
X2148 221 5 50 39 70 50 DFF_X1 $T=2330 12200 1 0 $X=2215 $Y=10685
X2149 183 5 50 39 174 50 DFF_X1 $T=2330 15000 1 0 $X=2215 $Y=13485
X2150 184 5 50 39 224 50 DFF_X1 $T=5560 6600 0 0 $X=5445 $Y=6485
X2151 197 9 50 39 225 50 DFF_X1 $T=12210 6600 0 0 $X=12095 $Y=6485
X2152 185 5 50 39 228 50 DFF_X1 $T=15440 6600 0 0 $X=15325 $Y=6485
X2153 186 5 50 39 124 50 DFF_X1 $T=18670 6600 0 0 $X=18555 $Y=6485
X2154 187 5 50 39 229 50 DFF_X1 $T=18670 9400 1 0 $X=18555 $Y=7885
X2155 198 9 50 39 126 50 DFF_X1 $T=22280 6600 0 0 $X=22165 $Y=6485
X2156 12 9 50 39 72 50 DFF_X1 $T=22280 9400 0 0 $X=22165 $Y=9285
X2210 114 1 50 39 363 50 AND2_X1 $T=1000 9400 1 0 $X=885 $Y=7885
X2211 114 2 50 39 313 50 AND2_X1 $T=1190 12200 1 0 $X=1075 $Y=10685
X2212 114 3 50 39 314 50 AND2_X1 $T=2330 9400 0 0 $X=2215 $Y=9285
X2213 67 222 50 39 340 50 AND2_X1 $T=6320 12200 0 0 $X=6205 $Y=12085
X2214 67 232 50 39 151 50 AND2_X1 $T=27790 6600 0 0 $X=27675 $Y=6485
X2215 95 260 50 39 261 50 AND2_X1 $T=55720 12200 1 0 $X=55605 $Y=10685
X2216 302 261 50 39 195 50 AND2_X1 $T=56670 9400 0 0 $X=56555 $Y=9285
X2217 105 369 50 39 104 50 AND2_X1 $T=63130 9400 0 180 $X=62255 $Y=7885
X2637 7 50 39 341 50 INV_X1 $T=7840 9400 1 0 $X=7725 $Y=7885
X2638 223 50 39 315 50 INV_X1 $T=9550 6600 0 0 $X=9435 $Y=6485
X2639 342 50 39 277 50 INV_X1 $T=10310 15000 1 0 $X=10195 $Y=13485
X2640 224 50 39 376 50 INV_X1 $T=10880 9400 1 0 $X=10765 $Y=7885
X2641 188 50 39 227 50 INV_X1 $T=11450 15000 1 0 $X=11335 $Y=13485
X2642 278 50 39 123 50 INV_X1 $T=11640 12200 0 0 $X=11525 $Y=12085
X2643 226 50 39 316 50 INV_X1 $T=12970 9400 1 0 $X=12855 $Y=7885
X2644 279 50 39 148 50 INV_X1 $T=14110 15000 1 0 $X=13995 $Y=13485
X2645 139 50 39 140 50 INV_X1 $T=14490 15000 1 0 $X=14375 $Y=13485
X2646 141 50 39 119 50 INV_X1 $T=15250 15000 0 180 $X=14755 $Y=13485
X2647 280 50 39 317 50 INV_X1 $T=20570 9400 0 0 $X=20455 $Y=9285
X2648 70 50 39 281 50 INV_X1 $T=23040 12200 1 0 $X=22925 $Y=10685
X2649 229 50 39 282 50 INV_X1 $T=23610 9400 1 0 $X=23495 $Y=7885
X2650 288 50 39 284 50 INV_X1 $T=24750 9400 1 0 $X=24635 $Y=7885
X2651 124 50 39 233 50 INV_X1 $T=25510 9400 1 0 $X=25395 $Y=7885
X2652 125 50 39 285 50 INV_X1 $T=25510 12200 0 0 $X=25395 $Y=12085
X2653 228 50 39 347 50 INV_X1 $T=25890 9400 1 0 $X=25775 $Y=7885
X2654 348 50 39 346 50 INV_X1 $T=26270 9400 1 0 $X=26155 $Y=7885
X2655 68 50 39 230 50 INV_X1 $T=26460 12200 0 0 $X=26345 $Y=12085
X2656 191 50 39 179 50 INV_X1 $T=28550 15000 0 180 $X=28055 $Y=13485
X2657 239 50 39 349 50 INV_X1 $T=30450 12200 0 0 $X=30335 $Y=12085
X2658 235 50 39 238 50 INV_X1 $T=30830 12200 0 0 $X=30715 $Y=12085
X2659 385 50 39 350 50 INV_X1 $T=32920 9400 0 0 $X=32805 $Y=9285
X2660 321 50 39 319 50 INV_X1 $T=34820 9400 0 0 $X=34705 $Y=9285
X2661 325 50 39 377 50 INV_X1 $T=44510 12200 1 180 $X=44015 $Y=12085
X2662 26 50 39 80 50 INV_X1 $T=46030 6600 1 180 $X=45535 $Y=6485
X2663 252 50 39 251 50 INV_X1 $T=46030 9400 1 0 $X=45915 $Y=7885
X2664 326 50 39 155 50 INV_X1 $T=46790 15000 0 180 $X=46295 $Y=13485
X2665 42 50 39 103 50 INV_X1 $T=47360 12200 1 180 $X=46865 $Y=12085
X2666 293 50 39 154 50 INV_X1 $T=47740 12200 1 180 $X=47245 $Y=12085
X2667 132 50 39 295 50 INV_X1 $T=48880 12200 1 180 $X=48385 $Y=12085
X2668 31 50 39 250 50 INV_X1 $T=49640 9400 1 0 $X=49525 $Y=7885
X2669 328 50 39 257 50 INV_X1 $T=50020 9400 0 0 $X=49905 $Y=9285
X2670 299 50 39 258 50 INV_X1 $T=52490 12200 0 180 $X=51995 $Y=10685
X2671 37 50 39 95 50 INV_X1 $T=54580 12200 0 0 $X=54465 $Y=12085
X2672 36 50 39 99 50 INV_X1 $T=54960 12200 0 0 $X=54845 $Y=12085
X2673 100 50 39 264 50 INV_X1 $T=58380 12200 0 0 $X=58265 $Y=12085
X2674 268 50 39 367 50 INV_X1 $T=60850 9400 1 0 $X=60735 $Y=7885
X2675 56 50 39 301 50 INV_X1 $T=61610 12200 0 180 $X=61115 $Y=10685
X2676 203 50 39 271 50 INV_X1 $T=61990 6600 1 180 $X=61495 $Y=6485
X2677 383 50 39 265 50 INV_X1 $T=64460 9400 1 180 $X=63965 $Y=9285
X2678 108 50 39 312 50 INV_X1 $T=64840 9400 0 180 $X=64345 $Y=7885
X2679 109 50 39 273 50 INV_X1 $T=65790 15000 0 180 $X=65295 $Y=13485
X2791 77 231 39 234 13 14 50 364 280 AOI222_X1 $T=28550 12200 1 0 $X=28435 $Y=10685
X2792 77 236 39 237 13 14 50 75 288 AOI222_X1 $T=31590 9400 0 180 $X=29955 $Y=7885
X2793 77 15 39 17 14 13 50 320 348 AOI222_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X2794 77 18 39 242 13 14 50 365 239 AOI222_X1 $T=34630 15000 0 180 $X=32995 $Y=13485
X2795 77 21 39 241 13 14 50 371 321 AOI222_X1 $T=33300 9400 0 0 $X=33185 $Y=9285
X2796 77 19 39 243 13 14 50 378 385 AOI222_X1 $T=38430 9400 0 0 $X=38315 $Y=9285
X2797 250 38 39 358 39 40 50 41 354 AOI222_X1 $T=53440 9400 1 0 $X=53325 $Y=7885
X2798 311 60 39 273 58 59 50 107 369 AOI222_X1 $T=62370 15000 1 0 $X=62255 $Y=13485
X2799 111 336 39 63 50 62 50 173 274 AOI222_X1 $T=67500 9400 0 180 $X=65865 $Y=7885
X2800 109 173 39 64 65 66 50 361 362 AOI222_X1 $T=66170 12200 0 0 $X=66055 $Y=12085
X2820 68 188 223 50 39 DLH_X1 $T=8980 12200 1 180 $X=6965 $Y=12085
X2821 68 342 7 50 39 DLH_X1 $T=7840 12200 1 0 $X=7725 $Y=10685
X2822 68 139 224 50 39 DLH_X1 $T=9740 12200 1 0 $X=9625 $Y=10685
X2823 68 278 8 50 39 DLH_X1 $T=11640 12200 1 0 $X=11525 $Y=10685
X2824 68 279 225 50 39 DLH_X1 $T=13540 12200 0 0 $X=13425 $Y=12085
X2825 68 143 226 50 39 DLH_X1 $T=13920 9400 0 0 $X=13805 $Y=9285
X2826 68 141 10 50 39 DLH_X1 $T=15820 12200 1 0 $X=15705 $Y=10685
X2827 68 190 11 50 39 DLH_X1 $T=20000 12200 0 0 $X=19885 $Y=12085
X2828 68 144 228 50 39 DLH_X1 $T=20570 12200 1 0 $X=20455 $Y=10685
X2829 68 145 229 50 39 DLH_X1 $T=22280 15000 1 0 $X=22165 $Y=13485
X2830 14 235 231 50 39 DLH_X1 $T=30450 15000 0 180 $X=28435 $Y=13485
X2831 14 16 236 50 39 DLH_X1 $T=31210 6600 1 180 $X=29195 $Y=6485
X2832 193 364 240 50 39 DLH_X1 $T=32540 12200 1 0 $X=32425 $Y=10685
X2833 14 26 20 50 39 DLH_X1 $T=39950 15000 0 180 $X=37935 $Y=13485
X2834 193 365 244 50 39 DLH_X1 $T=39380 12200 0 0 $X=39265 $Y=12085
X2835 14 55 19 50 39 DLH_X1 $T=39950 9400 1 0 $X=39835 $Y=7885
X2836 14 45 21 50 39 DLH_X1 $T=39950 9400 0 0 $X=39835 $Y=9285
X2837 14 29 18 50 39 DLH_X1 $T=39950 15000 1 0 $X=39835 $Y=13485
X2838 193 371 246 50 39 DLH_X1 $T=41850 9400 1 0 $X=41735 $Y=7885
X2839 193 378 248 50 39 DLH_X1 $T=43750 6600 0 0 $X=43635 $Y=6485
X2840 145 39 144 143 139 344 50 NOR4_X1 $T=17150 15000 0 180 $X=16085 $Y=13485
X2841 11 39 8 225 10 122 50 NOR4_X1 $T=18670 9400 1 180 $X=17605 $Y=9285
X2842 70 39 229 124 228 71 50 NOR4_X1 $T=24180 15000 1 0 $X=24065 $Y=13485
X2843 224 7 223 116 226 50 39 NOR4_X2 $T=10120 9400 0 0 $X=10005 $Y=9285
X2862 341 6 138 275 50 39 AOI21_X1 $T=8220 9400 1 0 $X=8105 $Y=7885
X2863 199 6 222 343 50 39 AOI21_X1 $T=8980 15000 1 0 $X=8865 $Y=13485
X2864 315 6 167 276 50 39 AOI21_X1 $T=9930 6600 0 0 $X=9815 $Y=6485
X2865 376 6 177 318 50 39 AOI21_X1 $T=12210 9400 1 0 $X=12095 $Y=7885
X2866 316 6 118 345 50 39 AOI21_X1 $T=13350 9400 1 0 $X=13235 $Y=7885
X2867 281 6 178 283 50 39 AOI21_X1 $T=23420 12200 1 0 $X=23305 $Y=10685
X2868 282 6 150 286 50 39 AOI21_X1 $T=23990 9400 1 0 $X=23875 $Y=7885
X2869 347 6 232 351 50 39 AOI21_X1 $T=26650 9400 1 0 $X=26535 $Y=7885
X2870 233 6 73 287 50 39 AOI21_X1 $T=28550 6600 0 0 $X=28435 $Y=6485
X2871 200 16 152 76 50 39 AOI21_X1 $T=33300 6600 0 0 $X=33185 $Y=6485
X2872 130 23 172 129 50 39 AOI21_X1 $T=42230 15000 1 0 $X=42115 $Y=13485
X2873 250 28 292 293 50 39 AOI21_X1 $T=46600 12200 1 0 $X=46485 $Y=10685
X2874 26 29 132 168 50 39 AOI21_X1 $T=46790 6600 0 0 $X=46675 $Y=6485
X2875 298 36 355 35 50 39 AOI21_X1 $T=51540 15000 1 0 $X=51425 $Y=13485
X2876 299 259 256 30 50 39 AOI21_X1 $T=53820 12200 0 0 $X=53705 $Y=12085
X2877 301 41 331 357 50 39 AOI21_X1 $T=55530 9400 1 180 $X=54655 $Y=9285
X2878 302 259 47 30 50 39 AOI21_X1 $T=57050 15000 1 0 $X=56935 $Y=13485
X2879 263 259 307 30 50 39 AOI21_X1 $T=58380 12200 1 180 $X=57505 $Y=12085
X2880 264 49 181 78 50 39 AOI21_X1 $T=58570 15000 0 180 $X=57695 $Y=13485
X2881 87 264 306 196 50 39 AOI21_X1 $T=59330 15000 0 180 $X=58455 $Y=13485
X2882 334 54 171 89 50 39 AOI21_X1 $T=60850 6600 1 180 $X=59975 $Y=6485
X2883 270 55 266 367 50 39 AOI21_X1 $T=61610 6600 1 180 $X=60735 $Y=6485
X2884 373 274 383 182 50 39 AOI21_X1 $T=65790 9400 1 180 $X=64915 $Y=9285
X2888 82 130 50 27 251 39 85 380 OAI221_X1 $T=46410 9400 1 0 $X=46295 $Y=7885
X2889 101 36 50 263 262 39 48 305 OAI221_X1 $T=58570 9400 1 180 $X=57315 $Y=9285
X2890 307 135 50 266 51 39 55 248 OAI221_X1 $T=58950 6600 0 0 $X=58835 $Y=6485
X2891 278 227 39 277 117 279 50 AOI22_X1 $T=11830 15000 1 0 $X=11715 $Y=13485
X2892 149 123 39 227 236 147 50 AOI22_X1 $T=20950 15000 0 180 $X=19885 $Y=13485
X2893 327 380 39 194 255 297 50 AOI22_X1 $T=47550 9400 1 0 $X=47435 $Y=7885
X2894 379 133 39 29 294 32 50 AOI22_X1 $T=49070 9400 0 0 $X=48955 $Y=9285
X2895 132 88 39 254 253 157 50 AOI22_X1 $T=49260 15000 1 0 $X=49145 $Y=13485
X2896 87 156 39 32 353 134 50 AOI22_X1 $T=49450 6600 0 0 $X=49335 $Y=6485
X2897 381 257 39 260 296 330 50 AOI22_X1 $T=50400 9400 0 0 $X=50285 $Y=9285
X2898 328 258 39 382 330 331 50 AOI22_X1 $T=51350 9400 0 0 $X=51235 $Y=9285
X2899 93 358 39 88 382 156 50 AOI22_X1 $T=54770 12200 1 0 $X=54655 $Y=10685
X2900 333 159 39 43 262 102 50 AOI22_X1 $T=57620 12200 1 0 $X=57505 $Y=10685
X2901 128 45 39 269 310 39 50 AOI22_X1 $T=62370 9400 0 0 $X=62255 $Y=9285
X2902 271 38 39 100 334 87 50 AOI22_X1 $T=65410 6600 1 180 $X=64345 $Y=6485
X2903 65 335 39 384 373 110 50 AOI22_X1 $T=67120 12200 0 180 $X=66055 $Y=10685
X2904 111 137 39 112 339 110 50 AOI22_X1 $T=69400 12200 1 180 $X=68335 $Y=12085
X2905 313 50 39 221 CLKBUF_X1 $T=1000 9400 0 0 $X=885 $Y=9285
X2906 363 50 39 375 CLKBUF_X1 $T=1380 6600 0 0 $X=1265 $Y=6485
X2907 314 50 39 374 CLKBUF_X1 $T=3660 9400 1 180 $X=2975 $Y=9285
X2908 69 120 50 343 230 142 39 OAI22_X1 $T=15250 15000 1 0 $X=15135 $Y=13485
X2909 69 225 50 275 230 317 39 OAI22_X1 $T=16770 9400 1 180 $X=15705 $Y=9285
X2910 69 8 50 276 230 284 39 OAI22_X1 $T=17720 9400 0 180 $X=16655 $Y=7885
X2911 69 10 50 318 230 285 39 OAI22_X1 $T=16770 9400 0 0 $X=16655 $Y=9285
X2912 69 11 50 345 230 346 39 OAI22_X1 $T=17720 9400 1 0 $X=17605 $Y=7885
X2913 147 148 50 231 277 149 39 OAI22_X1 $T=20950 15000 1 0 $X=20835 $Y=13485
X2914 69 126 50 286 230 349 39 OAI22_X1 $T=25510 12200 1 0 $X=25395 $Y=10685
X2915 69 72 50 283 230 205 39 OAI22_X1 $T=27220 15000 0 180 $X=26155 $Y=13485
X2916 69 192 50 351 230 350 39 OAI22_X1 $T=28360 9400 0 180 $X=27295 $Y=7885
X2917 69 74 50 287 230 319 39 OAI22_X1 $T=28740 9400 0 0 $X=28625 $Y=9285
X2918 78 80 50 290 130 82 39 OAI22_X1 $T=43940 9400 0 0 $X=43825 $Y=9285
X2919 136 361 50 311 57 56 39 OAI22_X1 $T=63320 12200 1 180 $X=62255 $Y=12085
X2930 290 29 39 245 247 50 202 291 AOI221_X1 $T=42230 12200 1 0 $X=42115 $Y=10685
X2931 250 98 39 35 257 50 170 368 AOI221_X1 $T=50970 9400 1 0 $X=50855 $Y=7885
X2932 258 35 39 37 368 50 300 357 AOI221_X1 $T=52300 9400 0 0 $X=52185 $Y=9285
X2933 42 55 39 46 35 50 49 263 AOI221_X1 $T=56480 12200 1 0 $X=56365 $Y=10685
X2934 337 107 39 61 39 50 269 165 AOI221_X1 $T=66170 12200 1 180 $X=64915 $Y=12085
X2935 76 238 240 352 50 39 50 OAI21_X1 $T=31780 12200 1 0 $X=31665 $Y=10685
X2936 292 252 379 103 50 39 50 OAI21_X1 $T=46600 9400 0 0 $X=46485 $Y=9285
X2937 131 30 324 295 50 39 50 OAI21_X1 $T=47740 12200 0 0 $X=47625 $Y=12085
X2938 329 34 297 256 50 39 50 OAI21_X1 $T=50780 12200 0 0 $X=50665 $Y=12085
X2939 148 50 342 175 39 NAND2_X1 $T=9740 15000 1 0 $X=9625 $Y=13485
X2940 279 50 277 176 39 NAND2_X1 $T=12590 12200 1 180 $X=11905 $Y=12085
X2941 76 50 238 352 39 NAND2_X1 $T=31780 12200 0 0 $X=31665 $Y=12085
X2942 79 50 84 83 39 NAND2_X1 $T=43750 15000 1 0 $X=43635 $Y=13485
X2943 25 50 84 293 39 NAND2_X1 $T=46790 15000 1 0 $X=46675 $Y=13485
X2944 294 50 45 327 39 NAND2_X1 $T=48120 6600 1 180 $X=47435 $Y=6485
X2945 80 50 23 169 39 NAND2_X1 $T=48500 6600 0 0 $X=48385 $Y=6485
X2946 253 50 86 249 39 NAND2_X1 $T=49260 15000 0 180 $X=48575 $Y=13485
X2947 295 50 50 298 39 NAND2_X1 $T=50210 12200 0 0 $X=50095 $Y=12085
X2948 355 50 158 254 39 NAND2_X1 $T=50780 15000 0 180 $X=50095 $Y=13485
X2949 257 50 33 329 39 NAND2_X1 $T=50780 12200 1 0 $X=50665 $Y=10685
X2950 90 50 45 356 39 NAND2_X1 $T=51730 6600 0 0 $X=51615 $Y=6485
X2951 96 50 91 92 39 NAND2_X1 $T=54010 15000 0 180 $X=53325 $Y=13485
X2952 101 50 32 360 39 NAND2_X1 $T=58570 9400 0 0 $X=58455 $Y=9285
X2953 128 50 27 332 39 NAND2_X1 $T=59710 12200 1 0 $X=59595 $Y=10685
X2954 272 50 103 309 39 NAND2_X1 $T=60850 12200 1 180 $X=60165 $Y=12085
X2955 50 50 166 338 39 NAND2_X1 $T=69020 15000 0 180 $X=68335 $Y=13485
X2956 83 39 28 260 50 NOR2_X1 $T=49260 12200 1 0 $X=49145 $Y=10685
X2957 46 39 27 299 50 NOR2_X1 $T=53060 12200 0 180 $X=52375 $Y=10685
X2958 34 39 94 259 50 NOR2_X1 $T=54010 15000 1 0 $X=53895 $Y=13485
X2959 46 39 35 42 50 302 NOR3_X1 $T=56100 12200 1 180 $X=55225 $Y=12085
X2960 50 127 207 352 39 XNOR2_X1 $T=31970 15000 1 0 $X=31855 $Y=13485
X2964 90 45 356 39 48 300 50 OAI211_X1 $T=52300 6600 0 0 $X=52185 $Y=6485
X2965 53 52 360 39 265 308 50 OAI211_X1 $T=60090 9400 1 180 $X=59025 $Y=9285
X2966 161 269 332 39 306 50 50 OAI211_X1 $T=61230 12200 0 180 $X=60165 $Y=10685
X2967 91 45 55 39 271 333 50 OAI211_X1 $T=61040 9400 0 0 $X=60925 $Y=9285
X2968 180 22 30 50 29 245 39 AOI211_X1 $T=41280 12200 0 0 $X=41165 $Y=12085
X2969 249 25 326 50 83 325 39 AOI211_X1 $T=46410 15000 0 180 $X=45345 $Y=13485
X2970 173 26 154 50 29 252 39 AOI211_X1 $T=45650 12200 1 0 $X=45535 $Y=10685
X2971 31 28 86 50 83 381 39 AOI211_X1 $T=49830 12200 1 0 $X=49715 $Y=10685
X2972 135 50 305 50 304 359 39 AOI211_X1 $T=58950 6600 1 180 $X=57885 $Y=6485
X2973 359 261 308 50 267 268 39 AOI211_X1 $T=61040 9400 1 180 $X=59975 $Y=9285
X2977 130 128 82 50 39 NOR2_X2 $T=40900 12200 1 0 $X=40785 $Y=10685
X2978 226 50 223 7 224 189 39 NAND4_X1 $T=10120 9400 1 180 $X=9055 $Y=9285
X2979 344 50 146 227 277 121 39 NAND4_X1 $T=17150 15000 1 0 $X=17035 $Y=13485
X2980 70 50 229 124 228 204 39 NAND4_X1 $T=24180 12200 0 0 $X=24065 $Y=12085
X2981 291 50 377 323 324 244 39 NAND4_X1 $T=43180 12200 0 0 $X=43065 $Y=12085
X2982 255 50 296 354 353 246 39 NAND4_X1 $T=50970 9400 0 180 $X=49905 $Y=7885
X2983 105 50 164 310 334 270 39 NAND4_X1 $T=63510 6600 0 0 $X=63395 $Y=6485
X2987 309 160 162 50 56 163 312 267 39 OAI33_X1 $T=60660 15000 1 0 $X=60545 $Y=13485
X2988 8 50 225 10 39 206 NAND3_X1 $T=18480 12200 0 180 $X=17605 $Y=10685
X2989 201 50 129 79 39 323 NAND3_X1 $T=42990 15000 1 0 $X=42875 $Y=13485
X2990 81 50 22 27 39 328 NAND3_X1 $T=44890 12200 1 0 $X=44775 $Y=10685
X2991 103 50 130 23 39 326 NAND3_X1 $T=46030 12200 1 180 $X=45155 $Y=12085
X2992 298 50 97 33 39 209 NAND3_X1 $T=51540 15000 0 180 $X=50665 $Y=13485
X2993 94 50 96 43 39 97 NAND3_X1 $T=55340 15000 1 0 $X=55225 $Y=13485
X2994 57 50 60 301 39 106 NAND3_X1 $T=63320 9400 0 0 $X=63205 $Y=9285
X2995 338 50 362 339 39 337 NAND3_X1 $T=68450 12200 1 180 $X=67575 $Y=12085
X3003 208 50 39 153 CLKBUF_X3 $T=42800 6600 0 0 $X=42685 $Y=6485
X3004 38 24 50 39 247 50 OR2_X1 $T=44130 12200 0 180 $X=43255 $Y=10685
X3005 234 370 231 50 39 191 50 HA_X1 $T=28740 12200 1 180 $X=26725 $Y=12085
X3006 237 372 236 50 39 370 50 HA_X1 $T=31590 9400 1 180 $X=29575 $Y=9285
X3007 241 366 21 50 39 289 50 HA_X1 $T=34440 12200 1 0 $X=34325 $Y=10685
X3008 320 322 15 50 39 372 50 HA_X1 $T=34630 9400 1 0 $X=34515 $Y=7885
X3009 242 20 18 50 39 366 50 HA_X1 $T=35200 12200 0 0 $X=35085 $Y=12085
X3010 243 289 19 50 39 322 50 HA_X1 $T=36720 6600 0 0 $X=36605 $Y=6485
X3011 358 29 45 50 39 269 50 HA_X1 $T=54960 9400 1 0 $X=54845 $Y=7885
X3012 272 269 55 50 39 361 50 HA_X1 $T=61610 12200 1 0 $X=61495 $Y=10685
X3013 336 271 55 50 39 137 50 HA_X1 $T=67120 6600 0 0 $X=67005 $Y=6485
X3014 335 100 55 50 39 64 50 HA_X1 $T=69020 12200 0 180 $X=67005 $Y=10685
X3015 384 45 55 50 39 112 50 HA_X1 $T=67500 9400 1 0 $X=67385 $Y=7885
.ENDS
***************************************
.SUBCKT CLKGATETST_X8 SE E CK GCK VSS VDD 7
** N=22 EP=7 IP=0 FDC=52
M0 8 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=170 $Y=90 $D=1
M1 VSS E 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=360 $Y=90 $D=1
M2 VSS 11 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=700 $Y=90 $D=1
M3 17 8 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=890 $Y=90 $D=1
M4 12 11 17 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.0125e-14 AS=3.85e-14 PD=8.7e-07 PS=8.3e-07 $X=1080 $Y=90 $D=1
M5 18 9 12 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.0125e-14 PD=4.6e-07 PS=8.7e-07 $X=1290 $Y=160 $D=1
M6 VSS 10 18 7 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=1480 $Y=160 $D=1
M7 10 12 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.58e-14 PD=1.11e-06 PS=1.12e-06 $X=1675 $Y=90 $D=1
M8 VSS 12 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1865 $Y=90 $D=1
M9 VSS CK 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=3.36e-14 PD=1.14e-06 PS=7.4e-07 $X=2260 $Y=90 $D=1
M10 19 CK VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=2465 $Y=90 $D=1
M11 13 12 19 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2655 $Y=90 $D=1
M12 20 12 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2845 $Y=90 $D=1
M13 VSS CK 20 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3035 $Y=90 $D=1
M14 21 CK VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3225 $Y=90 $D=1
M15 13 12 21 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3415 $Y=90 $D=1
M16 22 12 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3605 $Y=90 $D=1
M17 VSS CK 22 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=3795 $Y=90 $D=1
M18 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=3985 $Y=90 $D=1
M19 VSS 13 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4175 $Y=90 $D=1
M20 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4365 $Y=90 $D=1
M21 VSS 13 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4555 $Y=90 $D=1
M22 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4745 $Y=90 $D=1
M23 VSS 13 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=4935 $Y=90 $D=1
M24 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=5125 $Y=90 $D=1
M25 VSS 13 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=5315 $Y=90 $D=1
M26 14 SE 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=170 $Y=995 $D=0
M27 VDD E 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=360 $Y=995 $D=0
M28 VDD 11 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=700 $Y=995 $D=0
M29 15 8 VDD VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=890 $Y=890 $D=0
M30 12 9 15 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=4.245e-14 AS=5.88e-14 PD=1.16e-06 PS=1.12e-06 $X=1080 $Y=890 $D=0
M31 16 11 12 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=4.245e-14 PD=4.6e-07 PS=1.16e-06 $X=1290 $Y=1080 $D=0
M32 VDD 10 16 VDD PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=1480 $Y=1080 $D=0
M33 10 12 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=5.085e-14 PD=1.54e-06 PS=1.55e-06 $X=1675 $Y=680 $D=0
M34 VDD 12 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1865 $Y=680 $D=0
M35 VDD CK 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=5.04e-14 PD=1.57e-06 PS=9.5e-07 $X=2260 $Y=790 $D=0
M36 13 CK VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06 PS=1.57e-06 $X=2465 $Y=680 $D=0
M37 VDD 12 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2655 $Y=680 $D=0
M38 13 12 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2845 $Y=680 $D=0
M39 VDD CK 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3035 $Y=680 $D=0
M40 13 CK VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3225 $Y=680 $D=0
M41 VDD 12 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3415 $Y=680 $D=0
M42 13 12 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3605 $Y=680 $D=0
M43 VDD CK 13 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3795 $Y=680 $D=0
M44 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3985 $Y=680 $D=0
M45 VDD 13 GCK VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4175 $Y=680 $D=0
M46 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4365 $Y=680 $D=0
M47 VDD 13 GCK VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4555 $Y=680 $D=0
M48 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4745 $Y=680 $D=0
M49 VDD 13 GCK VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=4935 $Y=680 $D=0
M50 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=5125 $Y=680 $D=0
M51 VDD 13 GCK VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=5315 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125
** N=180 EP=124 IP=2370 FDC=1226
X1175 172 1 28 38 92 180 DFF_X1 $T=1000 1000 0 0 $X=885 $Y=885
X1176 168 2 28 38 79 28 DFF_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X1177 173 1 28 38 39 28 DFF_X1 $T=2330 3800 1 0 $X=2215 $Y=2285
X1178 174 1 28 38 93 180 DFF_X1 $T=8790 1000 0 0 $X=8675 $Y=885
X1179 152 9 28 38 41 28 DFF_X1 $T=9740 3800 0 0 $X=9625 $Y=3685
X1180 175 1 28 38 94 180 DFF_X1 $T=12020 1000 0 0 $X=11905 $Y=885
X1181 176 9 28 38 98 28 DFF_X1 $T=15440 3800 0 0 $X=15325 $Y=3685
X1182 126 9 28 38 44 28 DFF_X1 $T=18670 3800 1 0 $X=18555 $Y=2285
X1183 177 1 28 38 61 180 DFF_X1 $T=20380 1000 0 0 $X=20265 $Y=885
X1184 138 1 28 38 46 28 DFF_X1 $T=22280 3800 0 0 $X=22165 $Y=3685
X1185 139 9 28 38 100 28 DFF_X1 $T=25510 3800 0 0 $X=25395 $Y=3685
X1186 170 9 28 38 47 28 DFF_X1 $T=25890 6600 1 0 $X=25775 $Y=5085
X1187 103 1 28 38 95 180 DFF_X1 $T=27790 1000 0 0 $X=27675 $Y=885
X1188 169 1 28 38 108 180 DFF_X1 $T=34250 1000 1 180 $X=30905 $Y=885
X1189 104 1 28 38 96 28 DFF_X1 $T=36340 3800 0 0 $X=36225 $Y=3685
X1190 105 1 28 38 83 28 DFF_X1 $T=36720 6600 1 0 $X=36605 $Y=5085
X1191 118 1 28 38 63 180 DFF_X1 $T=40140 1000 1 180 $X=36795 $Y=885
X1274 60 3 28 38 151 28 AND2_X1 $T=3090 6600 0 180 $X=2215 $Y=5085
X1275 43 4 28 38 172 28 AND2_X1 $T=6130 3800 1 180 $X=5255 $Y=3685
X1276 60 5 28 38 157 28 AND2_X1 $T=6890 3800 1 180 $X=6015 $Y=3685
X1277 43 6 28 38 173 28 AND2_X1 $T=7650 3800 1 180 $X=6775 $Y=3685
X1278 43 7 28 38 174 28 AND2_X1 $T=7650 3800 0 0 $X=7535 $Y=3685
X1279 40 8 28 38 152 28 AND2_X1 $T=10690 3800 0 180 $X=9815 $Y=2285
X1280 40 10 28 38 42 28 AND2_X1 $T=12970 3800 1 0 $X=12855 $Y=2285
X1281 43 11 28 38 175 28 AND2_X1 $T=13730 3800 1 180 $X=12855 $Y=3685
X1282 40 12 28 38 176 180 AND2_X1 $T=16010 1000 1 180 $X=15135 $Y=885
X1283 40 13 28 38 126 180 AND2_X1 $T=17720 1000 0 0 $X=17605 $Y=885
X1284 60 14 28 38 137 28 AND2_X1 $T=19430 3800 1 180 $X=18555 $Y=3685
X1285 60 15 28 38 178 28 AND2_X1 $T=19430 3800 0 0 $X=19315 $Y=3685
X1286 60 16 28 38 158 28 AND2_X1 $T=19810 6600 1 0 $X=19695 $Y=5085
X1287 43 17 28 38 177 28 AND2_X1 $T=22660 6600 0 180 $X=21785 $Y=5085
X1288 43 18 28 38 138 28 AND2_X1 $T=22660 6600 1 0 $X=22545 $Y=5085
X1289 40 19 28 38 45 180 AND2_X1 $T=25320 1000 1 180 $X=24445 $Y=885
X1290 40 20 28 38 107 28 AND2_X1 $T=25130 6600 1 0 $X=25015 $Y=5085
X1291 40 21 28 38 139 180 AND2_X1 $T=25320 1000 0 0 $X=25205 $Y=885
X1292 40 22 28 38 170 180 AND2_X1 $T=27030 1000 0 0 $X=26915 $Y=885
X1293 40 23 28 38 80 28 AND2_X1 $T=30450 3800 0 0 $X=30335 $Y=3685
X1294 43 24 28 38 169 28 AND2_X1 $T=30640 6600 1 0 $X=30525 $Y=5085
X1295 40 25 28 38 62 28 AND2_X1 $T=33110 3800 1 0 $X=32995 $Y=2285
X1402 119 28 38 127 28 INV_X1 $T=34250 6600 0 180 $X=33755 $Y=5085
X1403 26 28 38 43 28 INV_X1 $T=39950 3800 1 180 $X=39455 $Y=3685
X1404 26 28 38 40 180 INV_X1 $T=40520 1000 1 180 $X=40025 $Y=885
X1405 30 28 38 49 28 INV_X1 $T=43750 6600 0 180 $X=43255 $Y=5085
X1406 140 28 38 128 28 INV_X1 $T=45270 3800 0 0 $X=45155 $Y=3685
X1407 37 28 38 29 180 INV_X1 $T=47550 1000 0 0 $X=47435 $Y=885
X1408 85 28 38 64 28 INV_X1 $T=50970 3800 1 0 $X=50855 $Y=2285
X1409 31 28 38 52 28 INV_X1 $T=51730 3800 1 0 $X=51615 $Y=2285
X1410 53 28 38 101 28 INV_X1 $T=53250 3800 1 180 $X=52755 $Y=3685
X1411 144 28 38 130 180 INV_X1 $T=54770 1000 1 180 $X=54275 $Y=885
X1412 71 28 38 34 28 INV_X1 $T=58000 3800 1 180 $X=57505 $Y=3685
X1413 147 28 38 135 28 INV_X1 $T=62370 3800 0 0 $X=62255 $Y=3685
X1414 155 28 38 134 180 INV_X1 $T=63700 1000 1 180 $X=63205 $Y=885
X1415 166 28 38 70 28 INV_X1 $T=63890 3800 1 0 $X=63775 $Y=2285
X1416 78 28 38 89 28 INV_X1 $T=64460 6600 0 180 $X=63965 $Y=5085
X1417 148 28 38 156 180 INV_X1 $T=65030 1000 0 0 $X=64915 $Y=885
X1469 109 81 127 28 38 DLH_X1 $T=32350 3800 0 0 $X=32235 $Y=3685
X1470 111 129 27 28 38 DLH_X1 $T=39950 6600 1 0 $X=39835 $Y=5085
X1471 109 112 128 28 38 DLH_X1 $T=41090 3800 0 0 $X=40975 $Y=3685
X1476 51 37 86 55 28 38 AOI21_X1 $T=51160 6600 1 0 $X=51045 $Y=5085
X1477 131 33 32 132 28 38 AOI21_X1 $T=53820 3800 0 0 $X=53705 $Y=3685
X1478 154 35 167 56 28 38 AOI21_X1 $T=60470 3800 0 0 $X=60355 $Y=3685
X1479 36 156 122 28 28 38 AOI21_X1 $T=61230 3800 0 0 $X=61115 $Y=3685
X1480 121 134 132 129 28 38 AOI21_X1 $T=62370 3800 1 0 $X=62255 $Y=2285
X1481 149 136 155 78 28 38 AOI21_X1 $T=64270 3800 1 0 $X=64155 $Y=2285
X1487 53 161 28 130 31 38 171 131 OAI221_X1 $T=53440 3800 1 0 $X=53325 $Y=2285
X1488 101 159 38 143 160 52 28 AOI22_X1 $T=51730 3800 0 0 $X=51615 $Y=3685
X1489 102 153 38 28 162 165 28 AOI22_X1 $T=56100 3800 0 180 $X=55035 $Y=2285
X1490 147 78 38 64 116 34 28 AOI22_X1 $T=58570 6600 1 0 $X=58455 $Y=5085
X1491 70 77 38 156 136 36 28 AOI22_X1 $T=65030 3800 1 0 $X=64915 $Y=2285
X1492 151 28 38 168 CLKBUF_X1 $T=3660 6600 0 180 $X=2975 $Y=5085
X1493 157 28 38 97 CLKBUF_X1 $T=4800 3800 0 0 $X=4685 $Y=3685
X1494 137 28 38 106 CLKBUF_X1 $T=19240 6600 0 180 $X=18555 $Y=5085
X1495 178 28 38 99 CLKBUF_X1 $T=20760 3800 1 180 $X=20075 $Y=3685
X1496 158 28 38 125 CLKBUF_X1 $T=21140 6600 0 180 $X=20455 $Y=5085
X1497 163 90 28 144 164 124 38 OAI22_X1 $T=57430 3800 1 0 $X=57315 $Y=2285
X1498 136 78 28 150 77 36 38 OAI22_X1 $T=66930 3800 0 180 $X=65865 $Y=2285
X1501 145 33 38 132 133 28 129 140 AOI221_X1 $T=55910 3800 0 0 $X=55795 $Y=3685
X1502 55 73 38 28 135 28 35 149 AOI221_X1 $T=62370 6600 1 0 $X=62255 $Y=5085
X1503 64 29 66 147 28 38 180 OAI21_X1 $T=47930 1000 0 0 $X=47815 $Y=885
X1504 28 30 87 85 28 38 28 OAI21_X1 $T=51920 6600 1 0 $X=51805 $Y=5085
X1505 70 89 115 146 28 38 28 OAI21_X1 $T=57620 6600 0 180 $X=56745 $Y=5085
X1506 70 28 69 147 38 NAND2_X1 $T=51730 3800 1 180 $X=51045 $Y=3685
X1507 160 28 162 145 38 NAND2_X1 $T=54580 3800 1 0 $X=54465 $Y=2285
X1508 29 28 89 71 38 NAND2_X1 $T=55340 6600 1 0 $X=55225 $Y=5085
X1509 55 28 89 114 38 NAND2_X1 $T=56480 6600 0 180 $X=55795 $Y=5085
X1510 34 28 49 146 38 NAND2_X1 $T=57620 3800 1 180 $X=56935 $Y=3685
X1511 34 28 64 154 38 NAND2_X1 $T=58760 3800 0 0 $X=58645 $Y=3685
X1512 49 28 29 166 38 NAND2_X1 $T=59520 3800 1 0 $X=59405 $Y=2285
X1513 36 28 148 74 38 NAND2_X1 $T=63510 6600 1 0 $X=63395 $Y=5085
X1514 32 38 82 110 28 NOR2_X1 $T=33300 6600 1 0 $X=33185 $Y=5085
X1515 51 38 37 55 28 NOR2_X1 $T=59520 6600 1 0 $X=59405 $Y=5085
X1516 26 60 28 38 INV_X2 $T=40140 3800 0 0 $X=40025 $Y=3685
X1519 150 28 76 167 75 133 38 NAND4_X1 $T=65220 3800 1 180 $X=64155 $Y=3685
X1533 48 26 28 38 141 180 OR2_X1 $T=41090 1000 0 0 $X=40975 $Y=885
X1534 48 26 28 38 179 28 OR2_X1 $T=41850 3800 0 180 $X=40975 $Y=2285
X1535 48 26 28 38 142 28 OR2_X1 $T=42230 3800 1 0 $X=42115 $Y=2285
X1536 120 84 30 28 38 51 28 HA_X1 $T=43750 6600 1 0 $X=43635 $Y=5085
X1537 159 114 129 28 38 161 180 HA_X1 $T=48690 1000 0 0 $X=48575 $Y=885
X1538 143 71 129 28 38 171 180 HA_X1 $T=52490 1000 0 0 $X=52375 $Y=885
X1539 72 85 37 28 38 88 28 HA_X1 $T=53440 6600 1 0 $X=53325 $Y=5085
X1540 153 146 129 28 38 164 180 HA_X1 $T=57050 1000 0 0 $X=56935 $Y=885
X1541 165 154 129 28 38 163 180 HA_X1 $T=58950 1000 0 0 $X=58835 $Y=885
X1542 54 51 37 28 38 148 180 HA_X1 $T=60850 1000 0 0 $X=60735 $Y=885
X1543 57 148 78 28 38 91 28 HA_X1 $T=64840 6600 1 0 $X=64725 $Y=5085
X1544 59 166 78 28 38 117 180 HA_X1 $T=67500 1000 0 0 $X=67385 $Y=885
X1545 123 147 78 28 38 58 28 HA_X1 $T=67500 3800 0 0 $X=67385 $Y=3685
X1546 28 141 65 67 28 38 28 CLKGATETST_X8 $T=45460 3800 1 0 $X=45345 $Y=2285
X1547 28 179 65 113 28 38 28 CLKGATETST_X8 $T=51160 3800 1 180 $X=45535 $Y=3685
X1548 28 142 65 68 28 38 28 CLKGATETST_X8 $T=45650 6600 1 0 $X=45535 $Y=5085
.ENDS
***************************************
.SUBCKT fpa_with_regisers VSS VDD inputB[18] inputB[17] inputA[18] inputB[16] inputA[17] inputA[16] inputB[15] inputB[0] inputB[9] inputA[15] inputB[11] inputA[9] inputB[8] inputB[10] inputA[10] inputA[8] inputB[2] inputB[3]
+ inputB[1] inputB[6] inputB[4] inputB[7] inputA[6] inputA[7] inputA[3] result[7] result[18] result[6] result[8] inputB[19] clk result[29] inputB[30] result[28] result[30] inputA[28] inputA[29] result[27]
+ inputA[30] inputB[26] inputA[27] inputB[25] inputB[24] result[24] result[23] inputA[26] inputA[25] inputA[24] inputA[23] result[26] inputA[14] result[25] inputA[12] result[13] result[12] result[14] en reset
+ result[2] result[16] result[4] result[17] result[3] result[1] result[5] inputA[5] result[10] inputA[2] result[9] inputA[4] inputA[11] result[11] result[0] inputA[0] inputB[5] result[15] inputA[1] inputA[13]
+ inputB[20] inputB[22] OF inputA[21] inputB[14] inputA[19] inputB[21] inputB[12] inputA[20] inputB[13] inputB[31] inputA[31] result[22] result[21] result[19] result[20] inputA[22] inputB[28] inputB[27] inputB[23]
+ result[31] inputB[29]
** N=732 EP=102 IP=1687 FDC=14720
X0 132 20 18 32 209 141 33 234 61 73 62 38 24 27 inputB[18] 34 42 200 29 41
+ inputB[17] 44 60 inputA[18] 52 120 75 inputB[16] 84 inputA[17] inputA[16] inputB[15] 76 74 80 inputB[0] 108 inputB[9] 104 78
+ inputA[15] 88 inputB[11] inputA[9] inputB[8] 89 92 inputA[10] 96 inputB[10] inputA[8] inputB[2] 91 inputB[1] inputB[7] inputB[3] inputB[4] inputB[6] inputA[6] 112
+ 114 inputA[7] 105 inputA[3] 687 14 VDD VSS 16 17 21 37 28 30 31 3 51 36 683 22
+ 39 143 43 123 64 285 69 97 115 119 result[6] result[3] 13 134 11 25 48 684 623 58
+ 68 86 99 81 result[4] result[17] 50 46 128 71 77 126 98 102 110 result[16] 53 56 65 70
+ 688 90 686 result[8] 26 59 127 result[18] result[7] result[2] 121 723 35 685 47 54 19 23 15 117
+ 624 12 66
+ ICV_8 $T=0 0 0 0 $X=0 $Y=59685
X1 132 22 18 136 139 34 144 38 143 60 71 140 724 33 26 690 27 4 175 138
+ 75 31 689 149 130 150 155 157 160 48 165 86 163 VSS 54 51 691 168 61 64
+ 90 62 69 162 102 181 304 631 176 167 81 74 84 76 693 98 196 183 187 92
+ 97 96 88 112 105 696 99 89 200 633 114 108 120 inputA[4] inputA[5] inputA[2] 687 2 VDD 21
+ 17 20 24 137 141 28 153 56 37 35 154 152 159 46 47 166 164 52 171 58
+ 184 66 65 173 174 73 179 177 80 129 186 191 192 194 195 199 119 123 135 209
+ 14 16 29 723 146 148 147 156 43 623 161 172 180 182 188 193 686 206 205 204
+ result[9] 133 13 11 142 25 12 145 185 53 697 197 208 131 44 685 169 695 190 624
+ result[10] result[5] 104 683 50 632 110 117 202 134 19 23 684 151 42 41 158 220 36 68
+ 170 121 result[1] 630 692 178 198 201 207 115 203 30 59 91 189 32 39 694 728
+ ICV_9 $T=0 0 0 0 $X=0 $Y=51260
X2 132 136 137 3 34 142 141 52 143 234 151 690 155 154 152 160 157 231 224 691
+ 168 5 236 56 64 167 181 226 304 252 2 228 631 298 239 170 81 171 73 242
+ 255 241 247 245 309 206 259 173 695 200 80 184 74 76 190 265 262 267 269 642
+ 696 257 192 189 inputB[5] 274 195 698 271 697 102 275 120 279 277 283 282 280 278 inputA[0]
+ inputA[1] inputA[11] 687 4 VSS VDD 11 17 135 140 212 24 138 18 144 147 689 148 150 221
+ 630 65 54 22 240 232 229 162 165 164 692 172 15 249 248 176 179 688 196 260
+ 272 264 266 198 203 202 201 119 123 209 724 134 217 29 149 146 218 225 156 254
+ 251 177 178 256 193 191 127 273 284 131 145 220 222 158 230 159 161 726 235 108
+ 244 243 246 180 694 188 197 285 268 result[11] result[15] 641 237 169 250 253 261 270 result[0] 133
+ 211 223 166 194 126 208 213 210 130 215 238 219 153 68 48 174 175 182 258 263
+ 633 281 139 227 163 729 78 632 186 199 70 185 187 693 204 205 207 183 276 214
+ 233
+ ICV_10 $T=0 0 0 0 $X=0 $Y=41485
X3 inputB[19] 200 287 120 inputA[13] 699 289 291 140 290 216 217 149 725 219 226 724 300 225 174
+ 4 141 130 224 181 304 308 303 231 298 228 223 52 307 54 311 238 700 317 315
+ 731 245 242 314 652 74 320 262 68 326 265 323 253 256 258 345 642 360 342 331
+ 330 423 338 267 703 365 269 332 363 364 VDD 270 701 343 195 702 429 698 8 352
+ 361 271 333 344 328 277 7 348 358 349 281 284 506 446 268 366 276 350 266 VSS
+ 285 214 138 145 295 689 150 222 301 179 144 229 240 569 128 172 243 80 76 247
+ 248 259 318 321 324 260 273 335 340 341 272 359 354 351 371 357 362 370 336 368
+ 279 210 132 211 123 288 213 3 218 220 299 221 155 227 29 230 237 316 263 261
+ 346 347 275 278 280 294 293 296 215 306 236 244 339 356 209 292 305 312 319 inputB[20]
+ 297 143 232 11 22 239 264 729 355 233 255 302 234 641 235 2 313 152 241 325
+ 327 129 334 353 283 212 250 329 322 251 337 369 249 246 252 257 274 367 310 282
+ 254 730
+ ICV_11 $T=0 0 0 0 $X=0 $Y=33085
X4 inputB[22] inputA[19] inputB[21] inputA[21] inputA[20] 200 120 inputB[13] inputB[14] 376 74 699 68 inputB[12] 289 288 375 380 140 391
+ 138 663 662 387 390 130 304 306 326 398 262 700 321 242 320 323 652 563 410 327
+ 413 417 325 359 666 330 408 418 331 704 421 422 358 506 430 424 708 266 348 709
+ 431 434 343 363 350 270 352 528 523 425 703 423 435 357 432 281 VSS 407 440 VDD
+ 344 342 429 441 442 443 447 362 366 284 8 346 351 349 285 373 80 290 378 295
+ 52 298 150 385 297 386 302 181 312 144 303 324 392 240 77 313 260 172 309 402
+ 394 404 319 328 412 416 702 401 333 706 405 707 337 335 339 414 340 426 338 341
+ 713 433 710 361 356 268 449 439 360 428 336 367 368 347 7 9 123 287 291 379
+ 294 381 296 217 384 382 229 388 389 305 307 329 492 409 334 345 711 354 364 365
+ 370 209 300 383 399 393 395 372 396 397 317 420 411 664 419 667 427 415 438 355
+ 445 369 374 400 665 437 444 448 299 728 314 705 292 226 179 318 332 353 224 228
+ 293 301 308 OF 406 403 273 687 712 311 322 446 377 315 310 701 436
+ ICV_12 $T=0 0 0 0 $X=0 $Y=24660
X5 inputB[31] inputA[31] 687 inputA[22] 120 373 375 74 456 716 376 68 454 460 461 470 475 479 482 485
+ 399 714 490 398 488 403 394 406 445 405 411 497 412 492 359 413 707 705 325 666
+ 501 415 410 327 428 503 422 708 432 338 436 505 VSS 513 510 425 348 270 370 523
+ 515 514 351 433 352 424 421 440 334 438 703 336 446 529 8 284 713 349 431 VDD
+ 119 465 459 463 662 468 18 386 304 472 389 474 160 476 174 396 727 316 715 481
+ 260 262 402 404 451 407 273 496 418 417 419 500 333 357 506 449 507 508 426 509
+ 342 511 528 347 518 512 521 581 430 276 710 439 331 719 437 328 711 363 356 441
+ 346 444 443 447 423 429 9 285 result[19] result[22] 374 457 458 381 466 383 464 382 290 384
+ 469 391 663 390 240 473 477 400 534 401 314 408 664 409 414 516 416 718 420 498
+ 706 665 504 427 434 268 435 522 266 525 712 531 123 result[21] 385 462 489 378 478 483
+ 484 315 487 326 330 493 494 495 519 343 709 524 675 732 455 139 480 499 717 502
+ 526 720 527 471 517 result[20] 80 379 388 5 393 486 704 533 448 453 467 297 387 395
+ 452 491 520 530 532 667 450 377 680 721 216 725 136 726 442 380 392
+ ICV_14 $T=0 0 0 0 $X=0 $Y=14840
X6 inputB[28] inputB[23] inputB[27] 687 200 74 537 543 120 542 476 549 262 326 471 556 558 489 473 490
+ 477 497 562 495 415 491 576 331 498 330 567 7 431 512 270 529 514 506 VDD 361
+ 575 407 363 578 585 519 371 521 527 VSS 583 357 577 580 591 440 722 362 532 526
+ 720 595 10 721 533 9 119 68 324 461 397 482 552 485 554 553 260 449 496 561
+ 499 492 718 421 702 513 343 423 511 572 370 680 522 276 515 516 517 570 581 590
+ 579 8 501 587 524 593 528 589 594 530 667 531 285 result[31] 730 716 541 463 465 382
+ 715 459 475 484 479 487 359 717 413 504 503 518 568 582 719 675 535 460 464 466
+ 467 468 472 474 470 174 462 304 550 551 557 560 507 502 573 508 338 681 523 336
+ 432 525 588 592 732 538 564 566 571 584 494 327 454 456 457 539 548 483 493 520
+ 428 453 536 544 545 546 458 727 469 486 481 273 565 574 350 540 547 455 555 500
+ 505 586 478 480 372 488 clk 510
+ ICV_15 $T=0 0 0 0 $X=0 $Y=6485
X7 687 200 inputB[29] 535 inputB[30] 538 539 inputA[28] 120 inputA[29] 541 inputA[30] inputA[27] inputB[26] inputB[25] inputB[24] 550 548 inputA[24] inputA[23]
+ inputA[26] inputA[25] inputA[14] 552 inputA[12] reset 471 VSS 576 498 517 555 574 580 279 361 585 VDD result[28] 123
+ 543 540 119 476 547 result[23] 485 en 562 578 571 680 575 586 584 589 594 10 285 result[24]
+ 450 result[14] 564 560 565 731 569 561 568 681 573 506 588 593 592 7 591 537 714 554
+ 556 result[12] 491 566 567 572 590 527 348 722 result[29] result[30] result[27] result[26] result[13] 536 542 545 481 570
+ 581 551 534 452 544 549 result[25] 273 553 326 558 563 577 579 582 732 451 557 505 587
+ 583 595 529 546
+ ICV_16 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
