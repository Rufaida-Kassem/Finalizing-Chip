* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SUPPLY_ERROR
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 9 A1 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 9 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q 6 7
** N=22 EP=7 IP=0 FDC=28
M0 VSS 11 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 19 10 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 9 8 19 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 20 11 9 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 20 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 10 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 21 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 12 8 21 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 22 11 12 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 14 22 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 14 12 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 12 QN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 14 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 11 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 15 10 VDD 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 9 11 15 7 PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 16 8 9 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 16 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 10 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 11 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 17 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 12 11 17 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 18 8 12 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 14 18 7 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 14 12 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 12 QN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 14 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5 6
** N=6 EP=6 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI222_X1 C2 C1 VDD B1 B2 A2 VSS A1 ZN 10 11
** N=16 EP=11 IP=0 FDC=12
M0 14 C2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN C1 14 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=1.2035e-13 AS=5.81e-14 PD=1.41e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 15 B1 ZN 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=1.2035e-13 PD=1.11e-06 PS=1.41e-06 $X=675 $Y=90 $D=1
M3 VSS B2 15 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=865 $Y=90 $D=1
M4 16 A2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1055 $Y=90 $D=1
M5 ZN A1 16 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1245 $Y=90 $D=1
M6 12 C2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD C1 12 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 12 B1 13 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=675 $Y=680 $D=0
M9 13 B2 12 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=865 $Y=680 $D=0
M10 ZN A2 13 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1055 $Y=680 $D=0
M11 13 A1 ZN 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1245 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT DLH_X1 G Q D VSS VDD 6 7
** N=15 EP=7 IP=0 FDC=16
M0 VSS G 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.205e-14 PD=1.11e-06 PS=6.3e-07 $X=170 $Y=90 $D=1
M1 Q 10 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS 8 9 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=755 $Y=215 $D=1
M3 14 D VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=945 $Y=215 $D=1
M4 10 9 14 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1135 $Y=215 $D=1
M5 15 8 10 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=1325 $Y=335 $D=1
M6 VSS 11 15 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=335 $D=1
M7 11 10 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=335 $D=1
M8 VDD G 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=170 $Y=995 $D=0
M9 Q 10 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M10 VDD 8 9 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=755 $Y=815 $D=0
M11 12 D VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=945 $Y=815 $D=0
M12 10 8 12 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1135 $Y=815 $D=0
M13 13 9 10 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=1325 $Y=1040 $D=0
M14 VDD 11 13 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=1.26e-14 PD=4.6e-07 PS=4.6e-07 $X=1515 $Y=1040 $D=0
M15 11 10 VDD 7 PMOS_VTL L=5e-08 W=9e-08 AD=9.45e-15 AS=1.26e-14 PD=3.9e-07 PS=4.6e-07 $X=1705 $Y=1040 $D=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 ZN A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 11 A3 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 10 A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 A3 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 12 A2 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 10 A2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI211_X1 C2 C1 A VDD B ZN VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 ZN C2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 10 C1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 12 A 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS B 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 11 C2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN C1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 VDD A ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 ZN B VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X3 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=8
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 7 Z 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=715 $Y=90 $D=1
M4 VDD A 7 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 VDD 7 Z 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN 8 9
** N=13 EP=9 IP=0 FDC=10
M0 10 A1 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 10 A3 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 10 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 A1 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 13 A3 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 13 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 10 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 10 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 9 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI22_X1 B2 B1 VDD A1 ZN A2 VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 11 B2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN B1 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 12 A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 VSS A2 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 VDD B2 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 10 B1 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 ZN A1 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 10 A2 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 VSS B2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 10 B1 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 10 A2 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 11 B2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 12 A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI221_X1 B2 B1 VSS A C2 VDD C1 ZN 9 10
** N=14 EP=10 IP=0 FDC=10
M0 VSS B2 11 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 B1 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 12 A 11 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN C2 12 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 12 C1 ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 13 B2 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 ZN B1 13 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 VDD A ZN 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 14 C2 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 ZN C1 14 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN B2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 9 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 10 B2 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6 7
** N=8 EP=7 IP=0 FDC=4
M0 8 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6 7
** N=8 EP=7 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 142
** N=247 EP=141 IP=3459 FDC=2148
X1475 65 1 58 57 201 241 244 AND2_X1 $T=1000 62600 1 0 $X=885 $Y=61085
X1476 76 143 58 57 203 242 245 AND2_X1 $T=6320 65400 1 180 $X=5445 $Y=65285
X1477 76 144 58 57 216 241 247 AND2_X1 $T=6130 62600 0 0 $X=6015 $Y=62485
X1478 76 145 58 57 231 242 245 AND2_X1 $T=7080 65400 1 180 $X=6205 $Y=65285
X1479 63 5 58 57 204 242 245 AND2_X1 $T=8220 65400 0 0 $X=8105 $Y=65285
X1480 76 146 58 57 207 242 245 AND2_X1 $T=10500 65400 0 0 $X=10385 $Y=65285
X1481 76 150 58 57 217 242 247 AND2_X1 $T=12780 65400 1 0 $X=12665 $Y=63885
X1482 65 12 58 57 151 243 245 AND2_X1 $T=13920 68200 0 180 $X=13045 $Y=66685
X1483 65 13 58 57 218 243 246 AND2_X1 $T=15820 68200 1 180 $X=14945 $Y=68085
X1484 65 15 58 57 219 243 246 AND2_X1 $T=16960 68200 0 0 $X=16845 $Y=68085
X1485 63 17 58 57 209 243 246 AND2_X1 $T=19620 68200 1 180 $X=18745 $Y=68085
X1486 63 18 58 57 233 243 246 AND2_X1 $T=20380 68200 1 180 $X=19505 $Y=68085
X1487 63 22 58 57 210 243 246 AND2_X1 $T=21900 68200 0 0 $X=21785 $Y=68085
X1488 65 26 58 57 220 243 246 AND2_X1 $T=27790 68200 1 180 $X=26915 $Y=68085
X1489 63 27 58 57 221 243 246 AND2_X1 $T=27790 68200 0 0 $X=27675 $Y=68085
X1490 65 29 58 57 211 243 246 AND2_X1 $T=29880 68200 0 0 $X=29765 $Y=68085
X1491 65 34 58 57 160 243 245 AND2_X1 $T=33490 68200 0 180 $X=32615 $Y=66685
X1492 65 37 58 57 162 243 246 AND2_X1 $T=33870 68200 0 0 $X=33755 $Y=68085
X1493 63 39 58 57 235 243 246 AND2_X1 $T=37290 68200 1 180 $X=36415 $Y=68085
X1494 63 41 58 57 189 243 246 AND2_X1 $T=38620 68200 0 0 $X=38505 $Y=68085
X1495 63 42 58 57 222 243 246 AND2_X1 $T=41660 68200 1 180 $X=40785 $Y=68085
X1496 63 43 58 57 191 243 246 AND2_X1 $T=41660 68200 0 0 $X=41545 $Y=68085
X1497 63 44 58 57 224 243 245 AND2_X1 $T=44320 68200 1 0 $X=44205 $Y=66685
X1498 65 45 58 57 223 243 246 AND2_X1 $T=44320 68200 0 0 $X=44205 $Y=68085
X1499 63 47 58 57 225 243 246 AND2_X1 $T=47550 68200 0 0 $X=47435 $Y=68085
X1500 65 103 58 57 226 243 246 AND2_X1 $T=50400 68200 1 180 $X=49525 $Y=68085
X1501 65 49 58 57 198 242 247 AND2_X1 $T=51920 65400 0 180 $X=51045 $Y=63885
X1502 65 50 58 57 212 243 246 AND2_X1 $T=51730 68200 0 0 $X=51615 $Y=68085
X1503 65 51 58 57 227 242 245 AND2_X1 $T=51920 65400 0 0 $X=51805 $Y=65285
X1504 65 52 58 57 193 242 247 AND2_X1 $T=54200 65400 0 180 $X=53325 $Y=63885
X1505 65 53 58 57 170 243 245 AND2_X1 $T=54580 68200 0 180 $X=53705 $Y=66685
X1506 63 54 58 57 228 243 246 AND2_X1 $T=57430 68200 1 180 $X=56555 $Y=68085
X1507 63 55 58 57 194 243 246 AND2_X1 $T=58950 68200 0 0 $X=58835 $Y=68085
X1508 76 200 58 57 215 242 245 AND2_X1 $T=59330 65400 0 0 $X=59215 $Y=65285
X1509 76 171 58 57 175 242 245 AND2_X1 $T=60090 65400 0 0 $X=59975 $Y=65285
X1510 76 172 58 57 229 241 247 AND2_X1 $T=62180 62600 1 180 $X=61305 $Y=62485
X1511 76 174 58 57 195 241 247 AND2_X1 $T=63890 62600 1 180 $X=63015 $Y=62485
X1512 76 173 58 57 199 242 247 AND2_X1 $T=63130 65400 1 0 $X=63015 $Y=63885
X1513 76 176 58 57 196 241 244 AND2_X1 $T=63890 62600 1 0 $X=63775 $Y=61085
X1514 76 177 58 57 230 241 247 AND2_X1 $T=63890 62600 0 0 $X=63775 $Y=62485
X1515 63 56 58 57 236 142 244 AND2_X1 $T=67120 59800 1 180 $X=66245 $Y=59685
X1527 201 3 58 57 152 241 247 DFF_X1 $T=1000 62600 0 0 $X=885 $Y=62485
X1528 216 4 58 57 113 242 245 DFF_X1 $T=1000 65400 0 0 $X=885 $Y=65285
X1529 203 4 58 57 128 243 245 DFF_X1 $T=1000 68200 1 0 $X=885 $Y=66685
X1530 231 4 58 57 114 243 245 DFF_X1 $T=7460 68200 0 180 $X=4115 $Y=66685
X1531 207 4 58 57 73 243 246 DFF_X1 $T=7270 68200 0 0 $X=7155 $Y=68085
X1532 204 7 58 57 16 242 247 DFF_X1 $T=7840 65400 1 0 $X=7725 $Y=63885
X1533 217 4 58 57 129 243 246 DFF_X1 $T=10500 68200 0 0 $X=10385 $Y=68085
X1534 151 3 58 57 153 242 245 DFF_X1 $T=14490 65400 1 180 $X=11145 $Y=65285
X1535 218 3 58 57 154 243 245 DFF_X1 $T=13920 68200 1 0 $X=13805 $Y=66685
X1536 219 3 58 57 155 242 245 DFF_X1 $T=14490 65400 0 0 $X=14375 $Y=65285
X1537 233 7 58 57 156 243 245 DFF_X1 $T=20380 68200 0 180 $X=17035 $Y=66685
X1538 209 7 58 57 24 242 247 DFF_X1 $T=21140 65400 1 0 $X=21025 $Y=63885
X1539 210 7 58 57 25 243 246 DFF_X1 $T=22660 68200 0 0 $X=22545 $Y=68085
X1540 220 3 58 57 158 242 245 DFF_X1 $T=24370 65400 0 0 $X=24255 $Y=65285
X1541 221 7 58 57 159 242 245 DFF_X1 $T=27600 65400 0 0 $X=27485 $Y=65285
X1542 160 3 58 57 161 242 247 DFF_X1 $T=30450 65400 1 0 $X=30335 $Y=63885
X1543 211 3 58 57 31 243 246 DFF_X1 $T=30640 68200 0 0 $X=30525 $Y=68085
X1544 235 7 58 57 96 243 245 DFF_X1 $T=36720 68200 0 180 $X=33375 $Y=66685
X1545 162 3 58 57 36 242 245 DFF_X1 $T=34250 65400 0 0 $X=34135 $Y=65285
X1546 222 7 58 57 166 243 245 DFF_X1 $T=36720 68200 1 0 $X=36605 $Y=66685
X1547 189 7 58 57 38 242 247 DFF_X1 $T=38050 65400 1 0 $X=37935 $Y=63885
X1548 191 7 58 57 167 242 247 DFF_X1 $T=41280 65400 1 0 $X=41165 $Y=63885
X1549 224 7 58 57 168 242 245 DFF_X1 $T=44700 65400 0 0 $X=44585 $Y=65285
X1550 223 3 58 57 163 243 245 DFF_X1 $T=45080 68200 1 0 $X=44965 $Y=66685
X1551 225 7 58 57 169 242 247 DFF_X1 $T=47930 65400 1 0 $X=47815 $Y=63885
X1552 226 3 58 57 164 243 245 DFF_X1 $T=48310 68200 1 0 $X=48195 $Y=66685
X1553 198 3 58 57 86 142 244 DFF_X1 $T=50400 59800 0 0 $X=50285 $Y=59685
X1554 227 3 58 57 28 241 247 DFF_X1 $T=50590 62600 0 0 $X=50475 $Y=62485
X1555 193 3 58 57 40 241 244 DFF_X1 $T=52490 62600 1 0 $X=52375 $Y=61085
X1556 212 3 58 57 165 243 246 DFF_X1 $T=52490 68200 0 0 $X=52375 $Y=68085
X1557 170 3 58 57 35 242 245 DFF_X1 $T=52680 65400 0 0 $X=52565 $Y=65285
X1558 199 4 58 57 110 241 244 DFF_X1 $T=60660 62600 0 180 $X=57315 $Y=61085
X1559 215 4 58 57 130 243 246 DFF_X1 $T=59710 68200 0 0 $X=59595 $Y=68085
X1560 228 7 58 57 81 242 247 DFF_X1 $T=59900 65400 1 0 $X=59785 $Y=63885
X1561 194 7 58 57 48 241 244 DFF_X1 $T=60660 62600 1 0 $X=60545 $Y=61085
X1562 229 4 58 57 111 242 245 DFF_X1 $T=62940 65400 0 0 $X=62825 $Y=65285
X1563 175 4 58 57 67 243 246 DFF_X1 $T=62940 68200 0 0 $X=62825 $Y=68085
X1564 236 7 58 57 87 142 244 DFF_X1 $T=66360 59800 1 180 $X=63015 $Y=59685
X1565 196 4 58 57 88 241 244 DFF_X1 $T=66170 62600 1 0 $X=66055 $Y=61085
X1566 195 4 58 57 101 241 247 DFF_X1 $T=66170 62600 0 0 $X=66055 $Y=62485
X1567 230 4 58 57 102 242 245 DFF_X1 $T=66170 65400 0 0 $X=66055 $Y=65285
X1768 152 58 57 183 241 247 INV_X1 $T=8220 62600 0 0 $X=8105 $Y=62485
X1769 206 58 57 143 241 247 INV_X1 $T=11070 62600 0 0 $X=10955 $Y=62485
X1770 186 58 57 145 242 247 INV_X1 $T=13540 65400 1 0 $X=13425 $Y=63885
X1771 208 58 57 146 241 247 INV_X1 $T=13730 62600 0 0 $X=13615 $Y=62485
X1772 179 58 57 150 242 247 INV_X1 $T=19240 65400 1 0 $X=19125 $Y=63885
X1773 108 58 57 188 142 244 INV_X1 $T=33110 59800 1 180 $X=32615 $Y=59685
X1774 238 58 57 200 242 245 INV_X1 $T=50780 65400 0 0 $X=50665 $Y=65285
X1775 239 58 57 171 241 247 INV_X1 $T=56480 62600 0 0 $X=56365 $Y=62485
X1776 237 58 57 173 241 247 INV_X1 $T=58380 62600 0 0 $X=58265 $Y=62485
X1777 213 58 57 172 241 247 INV_X1 $T=58760 62600 0 0 $X=58645 $Y=62485
X1778 214 58 57 174 142 244 INV_X1 $T=59140 59800 0 0 $X=59025 $Y=59685
X1779 240 58 57 176 142 244 INV_X1 $T=59520 59800 0 0 $X=59405 $Y=59685
X1780 140 58 57 177 142 244 INV_X1 $T=59900 59800 0 0 $X=59785 $Y=59685
X1795 112 156 57 6 154 19 58 135 206 241 247 AOI222_X1 $T=22280 62600 1 180 $X=20645 $Y=62485
X1796 112 24 57 6 155 19 58 64 208 241 244 AOI222_X1 $T=22660 62600 1 0 $X=22545 $Y=61085
X1797 112 25 57 6 153 19 58 136 186 241 247 AOI222_X1 $T=26460 62600 1 180 $X=24825 $Y=62485
X1798 112 159 57 6 158 19 58 137 179 241 247 AOI222_X1 $T=26460 62600 0 0 $X=26345 $Y=62485
X1799 112 167 57 6 161 46 58 132 238 241 247 AOI222_X1 $T=47550 62600 1 180 $X=45915 $Y=62485
X1800 112 166 57 6 31 46 58 138 239 241 247 AOI222_X1 $T=49070 62600 0 0 $X=48955 $Y=62485
X1801 112 168 57 6 163 46 58 100 213 241 244 AOI222_X1 $T=49450 62600 1 0 $X=49335 $Y=61085
X1802 112 169 57 6 164 46 58 85 237 241 244 AOI222_X1 $T=50970 62600 1 0 $X=50855 $Y=61085
X1803 112 48 57 6 165 46 58 139 214 142 244 AOI222_X1 $T=53630 59800 0 0 $X=53515 $Y=59685
X1804 112 81 57 6 35 46 58 66 240 142 244 AOI222_X1 $T=56670 59800 0 0 $X=56555 $Y=59685
X1823 19 91 152 58 57 241 247 DLH_X1 $T=14110 62600 0 0 $X=13995 $Y=62485
X1824 19 121 153 58 57 241 244 DLH_X1 $T=18100 62600 0 180 $X=16085 $Y=61085
X1825 19 78 16 58 57 142 244 DLH_X1 $T=17530 59800 0 0 $X=17415 $Y=59685
X1826 19 92 154 58 57 241 247 DLH_X1 $T=20760 62600 1 180 $X=18745 $Y=62485
X1827 19 122 155 58 57 241 244 DLH_X1 $T=20760 62600 1 0 $X=20645 $Y=61085
X1828 19 123 156 58 57 142 244 DLH_X1 $T=24560 59800 1 180 $X=22545 $Y=59685
X1829 19 106 158 58 57 241 244 DLH_X1 $T=27220 62600 1 0 $X=27105 $Y=61085
X1830 19 107 159 58 57 242 247 DLH_X1 $T=28550 65400 1 0 $X=28435 $Y=63885
X1831 19 72 28 58 57 241 244 DLH_X1 $T=29120 62600 1 0 $X=29005 $Y=61085
X1832 19 77 31 58 57 241 247 DLH_X1 $T=30640 62600 0 0 $X=30525 $Y=62485
X1833 46 125 161 58 57 241 247 DLH_X1 $T=32540 62600 0 0 $X=32425 $Y=62485
X1834 46 20 35 58 57 142 244 DLH_X1 $T=33110 59800 0 0 $X=32995 $Y=59685
X1835 46 108 36 58 57 241 244 DLH_X1 $T=33110 62600 1 0 $X=32995 $Y=61085
X1836 46 109 163 58 57 241 247 DLH_X1 $T=34440 62600 0 0 $X=34325 $Y=62485
X1837 46 33 38 58 57 241 244 DLH_X1 $T=35010 62600 1 0 $X=34895 $Y=61085
X1838 46 23 40 58 57 142 244 DLH_X1 $T=39000 59800 1 180 $X=36985 $Y=59685
X1839 46 79 164 58 57 241 244 DLH_X1 $T=38810 62600 1 0 $X=38695 $Y=61085
X1840 46 80 165 58 57 142 244 DLH_X1 $T=39000 59800 0 0 $X=38885 $Y=59685
X1841 46 97 166 58 57 241 247 DLH_X1 $T=42230 62600 1 180 $X=40215 $Y=62485
X1842 46 98 167 58 57 241 247 DLH_X1 $T=42230 62600 0 0 $X=42115 $Y=62485
X1843 46 99 168 58 57 142 244 DLH_X1 $T=45270 59800 1 180 $X=43255 $Y=59685
X1844 46 127 169 58 57 142 244 DLH_X1 $T=45270 59800 0 0 $X=45155 $Y=59685
X1845 46 84 48 58 57 142 244 DLH_X1 $T=48500 59800 0 0 $X=48385 $Y=59685
X1846 159 57 24 25 156 157 58 242 247 NOR4_X1 $T=26650 65400 0 180 $X=25585 $Y=63885
X1847 165 57 164 163 161 126 58 241 247 NOR4_X1 $T=39380 62600 0 0 $X=39265 $Y=62485
X1848 169 57 168 48 167 192 58 241 244 NOR4_X1 $T=46030 62600 1 0 $X=45915 $Y=61085
X1849 190 58 82 192 157 83 57 142 244 NAND4_X1 $T=42420 59800 0 0 $X=42305 $Y=59685
X1850 38 57 166 81 58 190 241 244 NOR3_X1 $T=41470 62600 1 0 $X=41355 $Y=61085
X1853 97 32 188 57 33 124 58 142 244 OAI211_X1 $T=31780 59800 0 0 $X=31665 $Y=59685
X1855 30 58 57 7 242 245 CLKBUF_X3 $T=31400 65400 0 0 $X=31285 $Y=65285
X1856 154 153 155 158 58 57 95 241 244 OR4_X1 $T=26080 62600 1 0 $X=25965 $Y=61085
X1857 133 2 180 202 58 57 142 244 AOI21_X1 $T=1760 59800 0 0 $X=1645 $Y=59685
X1858 70 2 197 89 58 57 142 244 AOI21_X1 $T=6890 59800 0 0 $X=6775 $Y=59685
X1859 183 6 144 116 58 57 241 247 AOI21_X1 $T=8600 62600 0 0 $X=8485 $Y=62485
X1860 187 14 131 232 58 57 241 244 AOI21_X1 $T=16200 62600 0 180 $X=15325 $Y=61085
X1861 21 20 93 185 58 57 142 244 AOI21_X1 $T=21900 59800 1 180 $X=21025 $Y=59685
X1862 21 23 94 234 58 57 142 244 AOI21_X1 $T=21900 59800 0 0 $X=21785 $Y=59685
X1864 180 68 57 69 205 104 58 142 244 AOI22_X1 $T=3090 59800 0 0 $X=2975 $Y=59685
X1865 115 68 57 69 184 180 58 241 244 AOI22_X1 $T=4610 62600 0 180 $X=3545 $Y=61085
X1866 115 69 57 68 149 181 58 241 244 AOI22_X1 $T=6130 62600 1 0 $X=6015 $Y=61085
X1867 197 71 57 69 62 59 58 142 244 AOI22_X1 $T=7650 59800 0 0 $X=7535 $Y=59685
X1868 59 68 57 69 187 181 58 241 244 AOI22_X1 $T=8790 62600 0 180 $X=7725 $Y=61085
X1869 205 14 57 72 147 21 58 142 244 AOI22_X1 $T=10690 59800 1 180 $X=9625 $Y=59685
X1870 9 105 57 14 148 184 58 241 244 AOI22_X1 $T=9930 62600 1 0 $X=9815 $Y=61085
X1871 117 14 57 105 118 11 58 142 244 AOI22_X1 $T=11830 59800 0 0 $X=11715 $Y=59685
X1872 60 105 57 14 178 149 58 241 247 AOI22_X1 $T=12400 62600 0 0 $X=12285 $Y=62485
X1873 90 105 57 14 119 62 58 142 244 AOI22_X1 $T=14300 59800 0 0 $X=14185 $Y=59685
X1874 61 105 57 77 120 21 58 142 244 AOI22_X1 $T=17530 59800 1 180 $X=16465 $Y=59685
X1875 61 75 58 232 10 187 57 241 244 OAI22_X1 $T=14490 62600 1 0 $X=14375 $Y=61085
X1876 205 10 58 147 8 57 72 74 142 244 OAI221_X1 $T=10690 59800 0 0 $X=10575 $Y=59685
X1877 184 10 58 148 9 57 75 234 241 244 OAI221_X1 $T=10880 62600 1 0 $X=10765 $Y=61085
X1878 60 75 58 178 149 57 10 185 241 244 OAI221_X1 $T=13160 62600 0 180 $X=11905 $Y=61085
X1880 70 2 181 182 58 57 241 244 OAI21_X1 $T=7080 62600 1 0 $X=6965 $Y=61085
X1881 134 58 2 182 57 142 244 NAND2_X1 $T=4990 59800 0 0 $X=4875 $Y=59685
X1882 134 57 2 202 58 142 244 NOR2_X1 $T=3090 59800 1 180 $X=2405 $Y=59685
.ENDS
***************************************
.SUBCKT ICV_7
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6 7
** N=11 EP=7 IP=0 FDC=10
M0 11 A 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 9 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 9 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 8 A VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 10 A ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 10 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8 9
** N=21 EP=9 IP=0 FDC=28
M0 VSS 10 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 19 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 10 A 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 11 CI 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 11 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 13 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 13 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 15 10 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 20 CI 15 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 21 B 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 21 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 15 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 10 CO 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 16 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 10 A 16 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 12 CI 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 12 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 14 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 14 A VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 15 10 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 17 CI 15 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 18 B 17 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 18 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 15 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI222_X1 C2 C1 VSS B1 B2 A2 VDD A1 ZN 10 11
** N=16 EP=11 IP=0 FDC=12
M0 12 C2 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS C1 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 12 B1 13 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=710 $Y=90 $D=1
M3 13 B2 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=900 $Y=90 $D=1
M4 ZN A2 13 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1090 $Y=90 $D=1
M5 13 A1 ZN 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1280 $Y=90 $D=1
M6 14 C2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M7 ZN C1 14 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M8 15 B1 ZN 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=710 $Y=680 $D=0
M9 VDD B2 15 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=900 $Y=680 $D=0
M10 16 A2 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1090 $Y=680 $D=0
M11 ZN A1 16 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1280 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN 9 10
** N=14 EP=10 IP=0 FDC=10
M0 13 B2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 13 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 14 C2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 14 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 11 B1 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 12 A 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 12 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 12 C1 ZN 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI211_X1 C2 C1 B VSS A ZN VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 12 C2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN C1 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS B ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN A VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 ZN C2 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 10 C1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 11 B 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=4
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 7 6 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 78 79 80 81
+ 82 83 84 85 86 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 211
+ 212
** N=369 EP=201 IP=4738 FDC=1742
X1852 117 251 73 72 280 366 369 AND2_X1 $T=52300 54200 0 0 $X=52185 $Y=54085
X1853 160 61 73 72 319 366 369 AND2_X1 $T=55720 54200 1 180 $X=54845 $Y=54085
X1854 117 254 73 72 321 365 369 AND2_X1 $T=63320 57000 1 0 $X=63205 $Y=55485
X1855 117 255 73 72 335 366 368 AND2_X1 $T=63510 54200 1 0 $X=63395 $Y=52685
X1856 117 256 73 72 322 211 367 AND2_X1 $T=63510 59800 1 0 $X=63395 $Y=58285
X1857 118 68 73 72 352 366 369 AND2_X1 $T=64080 54200 0 0 $X=63965 $Y=54085
X1858 118 69 73 72 353 366 368 AND2_X1 $T=64270 54200 1 0 $X=64155 $Y=52685
X1859 118 70 73 72 351 365 367 AND2_X1 $T=64460 57000 0 0 $X=64345 $Y=56885
X1874 319 59 73 72 237 365 369 DFF_X1 $T=56480 57000 0 180 $X=53135 $Y=55485
X1875 352 66 73 72 250 365 369 DFF_X1 $T=56480 57000 1 0 $X=56365 $Y=55485
X1876 353 66 73 72 249 366 369 DFF_X1 $T=58190 54200 0 0 $X=58075 $Y=54085
X1877 351 66 73 72 247 365 367 DFF_X1 $T=58190 57000 0 0 $X=58075 $Y=56885
X1878 335 71 73 72 179 212 368 DFF_X1 $T=66170 51400 0 0 $X=66055 $Y=51285
X1879 280 71 73 72 136 366 369 DFF_X1 $T=66170 54200 0 0 $X=66055 $Y=54085
X1880 321 71 73 72 119 365 369 DFF_X1 $T=66170 57000 1 0 $X=66055 $Y=55485
X1881 322 71 73 72 120 211 367 DFF_X1 $T=66170 59800 1 0 $X=66055 $Y=58285
X2305 199 73 72 338 366 369 INV_X1 $T=1380 54200 0 0 $X=1265 $Y=54085
X2306 2 73 72 3 366 368 INV_X1 $T=2520 54200 1 0 $X=2405 $Y=52685
X2307 257 73 72 122 365 369 INV_X1 $T=2900 57000 0 180 $X=2405 $Y=55485
X2308 289 73 72 285 211 367 INV_X1 $T=5180 59800 1 0 $X=5065 $Y=58285
X2309 262 73 72 213 366 369 INV_X1 $T=6890 54200 1 180 $X=6395 $Y=54085
X2310 291 73 72 181 211 367 INV_X1 $T=7270 59800 0 180 $X=6775 $Y=58285
X2311 292 73 72 290 365 369 INV_X1 $T=7460 57000 0 180 $X=6965 $Y=55485
X2312 294 73 72 325 366 368 INV_X1 $T=14490 54200 0 180 $X=13995 $Y=52685
X2313 189 73 72 104 212 368 INV_X1 $T=18480 51400 1 180 $X=17985 $Y=51285
X2314 298 73 72 267 366 368 INV_X1 $T=19050 54200 0 180 $X=18555 $Y=52685
X2315 303 73 72 297 365 369 INV_X1 $T=19240 57000 0 180 $X=18745 $Y=55485
X2316 299 73 72 344 366 368 INV_X1 $T=19810 54200 0 180 $X=19315 $Y=52685
X2317 300 73 72 327 211 367 INV_X1 $T=20190 59800 0 180 $X=19695 $Y=58285
X2318 150 73 72 343 212 368 INV_X1 $T=20380 51400 1 180 $X=19885 $Y=51285
X2319 302 73 72 222 212 368 INV_X1 $T=20760 51400 1 180 $X=20265 $Y=51285
X2320 78 73 72 306 365 367 INV_X1 $T=27410 57000 0 0 $X=27295 $Y=56885
X2321 83 73 72 174 212 368 INV_X1 $T=30640 51400 0 0 $X=30525 $Y=51285
X2322 24 73 72 84 211 367 INV_X1 $T=30830 59800 1 0 $X=30715 $Y=58285
X2323 191 73 72 184 212 368 INV_X1 $T=31020 51400 0 0 $X=30905 $Y=51285
X2324 217 73 72 358 366 368 INV_X1 $T=31020 54200 1 0 $X=30905 $Y=52685
X2325 192 73 72 175 212 368 INV_X1 $T=31400 51400 0 0 $X=31285 $Y=51285
X2326 34 73 72 231 365 367 INV_X1 $T=32920 57000 0 0 $X=32805 $Y=56885
X2327 215 73 72 276 366 368 INV_X1 $T=33680 54200 0 180 $X=33185 $Y=52685
X2328 110 73 72 235 365 369 INV_X1 $T=34440 57000 0 180 $X=33945 $Y=55485
X2329 228 73 72 307 211 367 INV_X1 $T=34630 59800 1 0 $X=34515 $Y=58285
X2330 227 73 72 229 365 369 INV_X1 $T=35390 57000 0 180 $X=34895 $Y=55485
X2331 12 73 72 274 211 367 INV_X1 $T=35010 59800 1 0 $X=34895 $Y=58285
X2332 48 73 72 233 366 368 INV_X1 $T=35200 54200 1 0 $X=35085 $Y=52685
X2333 47 73 72 277 366 368 INV_X1 $T=38050 54200 0 180 $X=37555 $Y=52685
X2334 112 73 72 185 211 367 INV_X1 $T=37860 59800 1 0 $X=37745 $Y=58285
X2335 29 73 72 278 212 368 INV_X1 $T=39190 51400 1 180 $X=38695 $Y=51285
X2336 51 73 72 330 365 367 INV_X1 $T=39570 57000 0 0 $X=39455 $Y=56885
X2337 193 73 72 239 211 367 INV_X1 $T=40140 59800 1 0 $X=40025 $Y=58285
X2338 317 73 72 316 366 368 INV_X1 $T=45080 54200 0 180 $X=44585 $Y=52685
X2339 157 73 72 86 366 369 INV_X1 $T=48310 54200 0 0 $X=48195 $Y=54085
X2340 195 73 72 158 366 369 INV_X1 $T=48690 54200 0 0 $X=48575 $Y=54085
X2341 318 73 72 159 365 369 INV_X1 $T=50970 57000 1 0 $X=50855 $Y=55485
X2342 196 73 72 186 366 369 INV_X1 $T=51920 54200 0 0 $X=51805 $Y=54085
X2343 197 73 72 336 366 369 INV_X1 $T=54960 54200 1 180 $X=54465 $Y=54085
X2344 91 73 72 178 365 367 INV_X1 $T=54770 57000 0 0 $X=54655 $Y=56885
X2345 334 73 72 350 366 369 INV_X1 $T=57430 54200 0 0 $X=57315 $Y=54085
X2346 198 73 72 282 366 369 INV_X1 $T=57810 54200 0 0 $X=57695 $Y=54085
X2347 253 73 72 92 365 367 INV_X1 $T=57810 57000 0 0 $X=57695 $Y=56885
X2348 281 73 72 254 365 369 INV_X1 $T=60090 57000 1 0 $X=59975 $Y=55485
X2349 320 73 72 256 211 367 INV_X1 $T=60090 59800 1 0 $X=59975 $Y=58285
X2350 283 73 72 255 366 368 INV_X1 $T=60470 54200 1 0 $X=60355 $Y=52685
X2403 9 215 72 4 6 7 73 124 214 366 368 AOI222_X1 $T=7460 54200 1 0 $X=7345 $Y=52685
X2404 9 110 72 10 6 7 73 75 216 366 369 AOI222_X1 $T=8600 54200 0 0 $X=8485 $Y=54085
X2405 7 13 72 12 9 6 73 8 324 365 367 AOI222_X1 $T=10310 57000 1 180 $X=8675 $Y=56885
X2406 9 217 72 11 6 7 73 97 262 366 368 AOI222_X1 $T=8980 54200 1 0 $X=8865 $Y=52685
X2407 7 137 72 14 6 9 73 24 292 365 369 AOI222_X1 $T=9930 57000 1 0 $X=9815 $Y=55485
X2408 9 15 72 138 6 7 73 165 364 365 367 AOI222_X1 $T=10310 57000 0 0 $X=10195 $Y=56885
X2409 41 226 72 140 31 32 73 172 225 212 368 AOI222_X1 $T=23990 51400 0 0 $X=23875 $Y=51285
X2410 41 227 72 33 31 32 73 80 223 366 369 AOI222_X1 $T=25890 54200 1 180 $X=24255 $Y=54085
X2411 41 236 72 37 31 32 73 182 361 366 369 AOI222_X1 $T=25890 54200 0 0 $X=25775 $Y=54085
X2412 41 228 72 38 31 32 73 183 329 212 368 AOI222_X1 $T=26460 51400 0 0 $X=26345 $Y=51285
X2413 32 46 72 40 41 31 73 153 268 366 369 AOI222_X1 $T=27410 54200 0 0 $X=27295 $Y=54085
X2414 32 188 72 42 31 41 73 49 224 366 368 AOI222_X1 $T=27790 54200 1 0 $X=27675 $Y=52685
X2415 308 363 72 45 46 47 73 278 201 212 368 AOI222_X1 $T=34820 51400 0 0 $X=34705 $Y=51285
X2416 90 54 72 248 55 56 73 88 318 212 368 AOI222_X1 $T=50020 51400 0 0 $X=49905 $Y=51285
X2417 60 247 72 58 39 53 73 336 320 365 367 AOI222_X1 $T=53250 57000 0 0 $X=53135 $Y=56885
X2418 60 249 72 58 237 53 73 135 283 366 368 AOI222_X1 $T=53630 54200 1 0 $X=53515 $Y=52685
X2419 90 248 72 62 55 56 73 252 253 366 368 AOI222_X1 $T=56670 54200 0 180 $X=55035 $Y=52685
X2420 60 250 72 58 63 53 73 350 281 365 367 AOI222_X1 $T=55150 57000 0 0 $X=55035 $Y=56885
X2421 60 57 72 58 64 53 73 282 93 211 367 AOI222_X1 $T=56670 59800 1 0 $X=56555 $Y=58285
X2422 90 62 72 65 55 56 73 187 334 212 368 AOI222_X1 $T=57050 51400 0 0 $X=56935 $Y=51285
X2468 151 80 30 73 72 365 369 DLH_X1 $T=23040 57000 1 0 $X=22925 $Y=55485
X2469 151 172 35 73 72 211 367 DLH_X1 $T=26650 59800 0 180 $X=24635 $Y=58285
X2470 151 217 39 73 72 211 367 DLH_X1 $T=26650 59800 1 0 $X=26535 $Y=58285
X2471 53 215 237 73 72 365 369 DLH_X1 $T=39950 57000 0 180 $X=37935 $Y=55485
X2472 53 228 52 73 72 211 367 DLH_X1 $T=40520 59800 1 0 $X=40405 $Y=58285
X2473 53 226 247 73 72 365 369 DLH_X1 $T=50970 57000 0 180 $X=48955 $Y=55485
X2474 53 48 249 73 72 366 368 DLH_X1 $T=50210 54200 1 0 $X=50095 $Y=52685
X2475 53 227 57 73 72 365 367 DLH_X1 $T=52300 57000 1 180 $X=50285 $Y=56885
X2476 53 236 250 73 72 365 369 DLH_X1 $T=51350 57000 1 0 $X=51235 $Y=55485
X2477 56 115 248 73 72 212 368 DLH_X1 $T=58570 51400 0 0 $X=58455 $Y=51285
X2478 116 252 67 73 72 212 368 DLH_X1 $T=60470 51400 0 0 $X=60355 $Y=51285
X2479 39 72 64 154 155 173 73 365 367 NOR4_X1 $T=27790 57000 0 0 $X=27675 $Y=56885
X2480 250 72 57 247 249 89 73 365 367 NOR4_X1 $T=52300 57000 0 0 $X=52185 $Y=56885
X2491 36 24 145 72 23 357 73 211 367 OAI211_X1 $T=17530 59800 0 180 $X=16465 $Y=58285
X2492 304 242 313 72 240 360 73 365 367 OAI211_X1 $T=40900 57000 1 180 $X=39835 $Y=56885
X2493 237 63 50 51 73 72 176 365 367 OR4_X1 $T=38430 57000 0 0 $X=38315 $Y=56885
X2494 285 1 180 323 73 72 211 367 AOI21_X1 $T=5560 59800 1 0 $X=5445 $Y=58285
X2495 325 19 293 166 73 72 212 368 AOI21_X1 $T=13920 51400 1 180 $X=13045 $Y=51285
X2496 344 22 356 127 73 72 366 369 AOI21_X1 $T=16770 54200 1 180 $X=15895 $Y=54085
X2497 222 22 342 301 73 72 365 369 AOI21_X1 $T=19240 57000 1 0 $X=19125 $Y=55485
X2498 28 29 305 340 73 72 366 369 AOI21_X1 $T=20760 54200 0 0 $X=20645 $Y=54085
X2499 269 22 303 328 73 72 365 369 AOI21_X1 $T=22280 57000 1 0 $X=22165 $Y=55485
X2500 28 215 271 270 73 72 365 367 AOI21_X1 $T=23040 57000 1 180 $X=22165 $Y=56885
X2501 28 15 346 355 73 72 211 367 AOI21_X1 $T=22280 59800 1 0 $X=22165 $Y=58285
X2502 28 217 272 362 73 72 365 367 AOI21_X1 $T=23040 57000 0 0 $X=22925 $Y=56885
X2503 236 231 349 359 73 72 365 369 AOI21_X1 $T=33490 57000 0 180 $X=32615 $Y=55485
X2504 360 243 133 314 73 72 366 369 AOI21_X1 $T=42990 54200 1 180 $X=42115 $Y=54085
X2506 121 2 72 3 94 337 73 212 368 AOI22_X1 $T=1000 51400 0 0 $X=885 $Y=51285
X2507 338 1 72 5 161 354 73 211 367 AOI22_X1 $T=1000 59800 1 0 $X=885 $Y=58285
X2508 354 1 72 5 95 285 73 211 367 AOI22_X1 $T=1950 59800 1 0 $X=1835 $Y=58285
X2509 122 5 72 1 259 258 73 365 367 AOI22_X1 $T=2140 57000 0 0 $X=2025 $Y=56885
X2510 123 1 72 5 260 258 73 212 368 AOI22_X1 $T=3470 51400 0 0 $X=3355 $Y=51285
X2511 161 96 72 74 18 259 73 211 367 AOI22_X1 $T=3850 59800 1 0 $X=3735 $Y=58285
X2512 259 96 72 74 264 288 73 365 369 AOI22_X1 $T=4230 57000 1 0 $X=4115 $Y=55485
X2513 260 96 72 74 287 142 73 212 368 AOI22_X1 $T=4420 51400 0 0 $X=4305 $Y=51285
X2514 261 2 72 3 162 216 73 365 367 AOI22_X1 $T=4420 57000 0 0 $X=4305 $Y=56885
X2515 260 74 72 96 221 288 73 366 368 AOI22_X1 $T=4610 54200 1 0 $X=4495 $Y=52685
X2516 164 3 72 2 289 143 73 212 368 AOI22_X1 $T=6320 51400 1 180 $X=5255 $Y=51285
X2517 163 2 72 3 257 214 73 366 368 AOI22_X1 $T=5560 54200 1 0 $X=5445 $Y=52685
X2518 7 14 72 137 337 9 73 366 368 AOI22_X1 $T=6510 54200 1 0 $X=6395 $Y=52685
X2519 214 2 72 3 291 324 73 365 367 AOI22_X1 $T=6700 57000 0 0 $X=6585 $Y=56885
X2520 7 138 72 165 261 9 73 365 369 AOI22_X1 $T=7460 57000 1 0 $X=7345 $Y=55485
X2521 125 98 72 100 218 287 73 212 368 AOI22_X1 $T=11070 51400 0 0 $X=10955 $Y=51285
X2522 263 98 72 100 219 221 73 366 368 AOI22_X1 $T=11830 54200 1 0 $X=11715 $Y=52685
X2523 264 100 72 98 220 265 73 365 369 AOI22_X1 $T=12590 57000 1 0 $X=12475 $Y=55485
X2524 342 103 72 101 167 341 73 365 367 AOI22_X1 $T=12970 57000 0 0 $X=12855 $Y=56885
X2525 295 103 72 101 168 266 73 366 369 AOI22_X1 $T=13160 54200 0 0 $X=13045 $Y=54085
X2526 341 103 72 101 294 295 73 366 368 AOI22_X1 $T=15440 54200 0 180 $X=14375 $Y=52685
X2527 126 101 72 103 263 144 73 212 368 AOI22_X1 $T=14680 51400 0 0 $X=14565 $Y=51285
X2528 266 103 72 101 265 144 73 366 369 AOI22_X1 $T=15060 54200 0 0 $X=14945 $Y=54085
X2529 104 22 72 27 266 343 73 212 368 AOI22_X1 $T=15630 51400 0 0 $X=15515 $Y=51285
X2530 326 103 72 101 169 342 73 365 367 AOI22_X1 $T=16960 57000 1 180 $X=15895 $Y=56885
X2531 356 296 72 101 20 297 73 365 369 AOI22_X1 $T=16390 57000 1 0 $X=16275 $Y=55485
X2532 343 22 72 27 341 267 73 366 368 AOI22_X1 $T=16770 54200 1 0 $X=16655 $Y=52685
X2533 267 22 72 27 326 344 73 366 369 AOI22_X1 $T=17720 54200 1 180 $X=16655 $Y=54085
X2534 326 101 72 103 170 297 73 365 367 AOI22_X1 $T=16960 57000 0 0 $X=16845 $Y=56885
X2535 171 22 72 27 295 222 73 366 368 AOI22_X1 $T=17720 54200 1 0 $X=17605 $Y=52685
X2536 223 106 72 107 298 105 73 366 368 AOI22_X1 $T=20760 54200 0 180 $X=19695 $Y=52685
X2537 78 147 72 26 300 306 73 365 367 AOI22_X1 $T=21140 57000 1 180 $X=20075 $Y=56885
X2538 129 107 72 106 302 225 73 212 368 AOI22_X1 $T=22090 51400 0 0 $X=21975 $Y=51285
X2539 361 106 72 107 269 79 73 366 368 AOI22_X1 $T=22850 54200 1 0 $X=22735 $Y=52685
X2540 329 106 72 107 299 152 73 212 368 AOI22_X1 $T=23040 51400 0 0 $X=22925 $Y=51285
X2541 32 153 72 46 105 41 73 212 368 AOI22_X1 $T=25510 51400 0 0 $X=25395 $Y=51285
X2542 131 15 72 40 275 306 73 365 369 AOI22_X1 $T=30260 57000 1 0 $X=30145 $Y=55485
X2543 131 24 72 49 347 306 73 365 367 AOI22_X1 $T=30260 57000 0 0 $X=30145 $Y=56885
X2544 131 34 72 236 279 306 73 366 369 AOI22_X1 $T=30450 54200 0 0 $X=30335 $Y=54085
X2545 131 217 72 226 273 306 73 366 369 AOI22_X1 $T=31400 54200 0 0 $X=31285 $Y=54085
X2546 49 84 72 274 348 228 73 211 367 AOI22_X1 $T=31780 59800 1 0 $X=31665 $Y=58285
X2547 48 276 72 358 230 226 73 366 368 AOI22_X1 $T=32350 54200 1 0 $X=32235 $Y=52685
X2548 348 109 72 12 359 307 73 211 367 AOI22_X1 $T=32730 59800 1 0 $X=32615 $Y=58285
X2549 304 242 72 345 243 315 73 365 369 AOI22_X1 $T=41280 57000 1 0 $X=41165 $Y=55485
X2550 245 309 72 82 156 114 73 366 368 AOI22_X1 $T=41850 54200 1 0 $X=41735 $Y=52685
X2551 55 54 72 85 317 90 73 212 368 AOI22_X1 $T=50020 51400 1 180 $X=48955 $Y=51285
X2552 25 146 73 148 149 327 72 365 367 OAI22_X1 $T=19240 57000 0 0 $X=19125 $Y=56885
X2553 227 235 73 232 231 236 72 366 369 OAI22_X1 $T=34440 54200 1 180 $X=33375 $Y=54085
X2554 245 309 73 241 312 311 72 366 368 OAI22_X1 $T=40900 54200 0 180 $X=39835 $Y=52685
X2555 364 2 73 5 216 72 3 200 365 367 OAI221_X1 $T=8790 57000 1 180 $X=7535 $Y=56885
X2556 264 102 73 220 265 72 16 270 365 367 OAI221_X1 $T=12970 57000 1 180 $X=11715 $Y=56885
X2557 125 16 73 218 287 72 102 99 212 368 OAI221_X1 $T=12020 51400 0 0 $X=11905 $Y=51285
X2558 263 16 73 219 221 72 102 340 366 369 OAI221_X1 $T=12020 54200 0 0 $X=11905 $Y=54085
X2559 168 16 73 17 18 72 102 362 211 367 OAI221_X1 $T=12590 59800 1 0 $X=12475 $Y=58285
X2560 76 102 73 21 20 72 16 355 211 367 OAI221_X1 $T=14870 59800 0 180 $X=13615 $Y=58285
X2561 268 107 73 27 223 72 106 296 366 369 OAI221_X1 $T=19620 54200 0 0 $X=19505 $Y=54085
X2562 232 349 73 230 229 72 110 363 366 369 OAI221_X1 $T=33490 54200 1 180 $X=32235 $Y=54085
X2563 330 113 73 238 239 72 25 251 366 368 OAI221_X1 $T=38810 54200 1 0 $X=38695 $Y=52685
X2565 338 1 288 339 73 72 366 369 OAI21_X1 $T=1760 54200 0 0 $X=1645 $Y=54085
X2566 213 2 354 284 73 72 365 369 OAI21_X1 $T=1760 57000 1 0 $X=1645 $Y=55485
X2567 141 3 258 286 73 72 366 369 OAI21_X1 $T=3090 54200 0 0 $X=2975 $Y=54085
X2568 325 139 245 293 73 72 212 368 OAI21_X1 $T=13920 51400 0 0 $X=13805 $Y=51285
X2569 36 12 304 108 73 72 211 367 OAI21_X1 $T=23990 59800 1 0 $X=23875 $Y=58285
X2570 36 34 345 81 73 72 365 367 OAI21_X1 $T=26080 57000 1 180 $X=25205 $Y=56885
X2571 36 15 313 346 73 72 365 367 OAI21_X1 $T=26080 57000 0 0 $X=25965 $Y=56885
X2572 36 215 82 271 73 72 365 369 OAI21_X1 $T=27600 57000 0 180 $X=26725 $Y=55485
X2573 36 217 312 272 73 72 365 369 OAI21_X1 $T=27600 57000 1 0 $X=27485 $Y=55485
X2574 36 29 130 305 73 72 366 368 OAI21_X1 $T=29310 54200 1 0 $X=29195 $Y=52685
X2575 44 40 240 275 73 72 365 369 OAI21_X1 $T=35390 57000 1 0 $X=35275 $Y=55485
X2576 44 236 315 279 73 72 366 369 OAI21_X1 $T=37100 54200 0 0 $X=36985 $Y=54085
X2577 44 49 310 347 73 72 365 367 OAI21_X1 $T=37670 57000 0 0 $X=37555 $Y=56885
X2578 44 226 311 273 73 72 366 368 OAI21_X1 $T=38050 54200 1 0 $X=37935 $Y=52685
X2579 94 73 1 339 72 366 368 NAND2_X1 $T=1950 54200 1 0 $X=1835 $Y=52685
X2580 337 73 2 284 72 366 369 NAND2_X1 $T=3090 54200 1 180 $X=2405 $Y=54085
X2581 261 73 3 286 72 366 369 NAND2_X1 $T=4420 54200 1 180 $X=3735 $Y=54085
X2582 316 73 53 238 72 366 368 NAND2_X1 $T=43370 54200 0 180 $X=42685 $Y=52685
X2583 269 72 22 301 73 365 369 NOR2_X1 $T=21140 57000 0 180 $X=20455 $Y=55485
X2584 241 72 194 132 73 212 368 NOR2_X1 $T=40900 51400 0 0 $X=40785 $Y=51285
X2585 315 72 345 314 73 366 369 NOR2_X1 $T=42230 54200 1 180 $X=41545 $Y=54085
X2603 73 147 128 26 72 211 367 XNOR2_X1 $T=19810 59800 0 180 $X=18555 $Y=58285
X2604 73 315 333 332 72 366 369 XNOR2_X1 $T=44130 54200 0 0 $X=44015 $Y=54085
X2605 73 345 62 333 72 366 369 XNOR2_X1 $T=48310 54200 1 180 $X=47055 $Y=54085
X2606 331 244 310 357 72 73 54 365 367 FA_X1 $T=43940 57000 1 180 $X=40785 $Y=56885
X2607 246 245 309 133 72 73 65 212 368 FA_X1 $T=44510 51400 1 180 $X=41355 $Y=51285
X2608 332 331 242 304 72 73 248 365 369 FA_X1 $T=45270 57000 0 180 $X=42115 $Y=55485
X2609 244 313 240 73 72 73 85 365 367 FA_X1 $T=43940 57000 0 0 $X=43825 $Y=56885
X2610 134 246 311 312 72 73 177 366 368 FA_X1 $T=48120 54200 0 180 $X=44965 $Y=52685
X2617 78 229 73 227 44 43 72 235 309 366 369 OAI222_X1 $T=35960 54200 1 180 $X=34325 $Y=54085
X2618 78 307 73 228 44 43 72 274 242 365 367 OAI222_X1 $T=34820 57000 0 0 $X=34705 $Y=56885
X2619 78 233 73 48 44 43 72 276 114 366 368 OAI222_X1 $T=35580 54200 1 0 $X=35465 $Y=52685
X2620 78 277 73 47 44 43 72 278 111 212 368 OAI222_X1 $T=36340 51400 0 0 $X=36225 $Y=51285
X2623 290 3 72 1 213 73 2 323 365 369 AOI221_X1 $T=5180 57000 1 0 $X=5065 $Y=55485
X2624 224 106 72 22 225 73 107 328 366 369 AOI221_X1 $T=21520 54200 0 0 $X=21405 $Y=54085
X2625 277 29 72 234 233 73 215 308 366 368 AOI221_X1 $T=34820 54200 0 180 $X=33565 $Y=52685
X2626 48 276 226 73 358 234 72 212 368 AOI211_X1 $T=32160 51400 0 0 $X=32045 $Y=51285
X2627 190 73 72 151 365 367 CLKBUF_X1 $T=29500 57000 0 0 $X=29385 $Y=56885
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X2 A ZN VSS VDD 5 6
** N=6 EP=6 IP=0 FDC=4
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A ZN 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A ZN 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI33_X1 B3 B2 B1 VSS A1 A2 A3 ZN VDD 10 11
** N=16 EP=11 IP=0 FDC=12
M0 12 B3 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS B2 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 12 B1 VSS 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 ZN A1 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 12 A2 ZN 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 ZN A3 12 10 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1110 $Y=90 $D=1
M6 13 B3 VDD 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M7 14 B2 13 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M8 ZN B1 14 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M9 15 A1 ZN 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M10 16 A2 15 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
M11 VDD A3 16 11 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1110 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X2 A1 ZN A2 VSS VDD 6 7
** N=9 EP=7 IP=0 FDC=8
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 ZN A1 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 VSS A2 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=755 $Y=90 $D=1
M4 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M5 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M6 9 A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M7 VDD A2 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=755 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202
+ 223 224
** N=368 EP=202 IP=4779 FDC=1824
X1916 90 268 68 67 356 364 366 AND2_X1 $T=60470 45800 0 0 $X=60355 $Y=45685
X1917 153 58 68 67 270 364 366 AND2_X1 $T=63130 45800 0 0 $X=63015 $Y=45685
X1918 90 269 68 67 357 365 367 AND2_X1 $T=63320 48600 0 0 $X=63205 $Y=48485
X1919 116 64 68 67 271 364 368 AND2_X1 $T=66550 45800 1 0 $X=66435 $Y=44285
X1932 162 45 68 67 126 223 368 DFF_X1 $T=42420 43000 0 0 $X=42305 $Y=42885
X1933 271 65 68 67 160 223 368 DFF_X1 $T=66170 43000 0 0 $X=66055 $Y=42885
X1934 163 66 68 67 161 364 366 DFF_X1 $T=66170 45800 0 0 $X=66055 $Y=45685
X1935 356 66 68 67 181 365 366 DFF_X1 $T=66170 48600 1 0 $X=66055 $Y=47085
X1936 357 66 68 67 117 224 367 DFF_X1 $T=66170 51400 1 0 $X=66055 $Y=49885
X2369 358 68 67 330 365 367 INV_X1 $T=1760 48600 0 0 $X=1645 $Y=48485
X2370 300 68 67 274 223 368 INV_X1 $T=2710 43000 0 0 $X=2595 $Y=42885
X2371 139 68 67 138 224 367 INV_X1 $T=3850 51400 0 180 $X=3355 $Y=49885
X2372 307 68 67 70 365 367 INV_X1 $T=6700 48600 1 180 $X=6205 $Y=48485
X2373 75 68 67 13 223 368 INV_X1 $T=17910 43000 0 0 $X=17795 $Y=42885
X2374 315 68 67 100 224 367 INV_X1 $T=19620 51400 0 180 $X=19125 $Y=49885
X2375 17 68 67 77 364 366 INV_X1 $T=22660 45800 1 180 $X=22165 $Y=45685
X2376 123 68 67 26 223 368 INV_X1 $T=24560 43000 0 0 $X=24445 $Y=42885
X2377 12 68 67 239 364 368 INV_X1 $T=25510 45800 1 0 $X=25395 $Y=44285
X2378 78 68 67 287 364 368 INV_X1 $T=25890 45800 1 0 $X=25775 $Y=44285
X2379 31 68 67 318 365 367 INV_X1 $T=26840 48600 0 0 $X=26725 $Y=48485
X2380 14 68 67 238 364 366 INV_X1 $T=27790 45800 1 180 $X=27295 $Y=45685
X2381 33 68 67 322 365 366 INV_X1 $T=31020 48600 0 180 $X=30525 $Y=47085
X2382 15 68 67 244 365 367 INV_X1 $T=31020 48600 1 180 $X=30525 $Y=48485
X2383 351 68 67 360 224 367 INV_X1 $T=32730 51400 0 180 $X=32235 $Y=49885
X2384 35 68 67 290 365 367 INV_X1 $T=32540 48600 0 0 $X=32425 $Y=48485
X2385 11 68 67 248 365 367 INV_X1 $T=33300 48600 1 180 $X=32805 $Y=48485
X2386 3 68 67 247 365 367 INV_X1 $T=33300 48600 0 0 $X=33185 $Y=48485
X2387 36 68 67 251 365 367 INV_X1 $T=35580 48600 1 180 $X=35085 $Y=48485
X2388 291 68 67 353 364 368 INV_X1 $T=37860 45800 0 180 $X=37365 $Y=44285
X2389 38 68 67 252 365 367 INV_X1 $T=37670 48600 0 0 $X=37555 $Y=48485
X2390 16 68 67 39 224 367 INV_X1 $T=39570 51400 0 180 $X=39075 $Y=49885
X2391 355 68 67 292 365 367 INV_X1 $T=42420 48600 1 180 $X=41925 $Y=48485
X2392 86 68 67 268 364 368 INV_X1 $T=50400 45800 1 0 $X=50285 $Y=44285
X2393 194 68 67 269 364 366 INV_X1 $T=54010 45800 0 0 $X=53895 $Y=45685
X2394 298 68 67 187 224 367 INV_X1 $T=54580 51400 1 0 $X=54465 $Y=49885
X2457 5 9 67 132 6 74 68 4 120 364 366 AOI222_X1 $T=9550 45800 1 180 $X=7915 $Y=45685
X2458 5 7 67 8 6 74 68 15 182 224 367 AOI222_X1 $T=8220 51400 1 0 $X=8105 $Y=49885
X2459 25 19 67 20 21 22 68 23 171 364 366 AOI222_X1 $T=22660 45800 0 0 $X=22545 $Y=45685
X2460 21 133 67 24 22 25 68 123 184 224 367 AOI222_X1 $T=24180 51400 1 0 $X=24065 $Y=49885
X2461 87 44 67 40 41 43 68 192 196 223 368 AOI222_X1 $T=40900 43000 0 0 $X=40785 $Y=42885
X2462 87 260 67 44 41 43 68 125 85 364 368 AOI222_X1 $T=42610 45800 1 0 $X=42495 $Y=44285
X2463 87 261 67 260 41 43 68 296 197 364 368 AOI222_X1 $T=46030 45800 1 0 $X=45915 $Y=44285
X2464 87 263 67 261 41 43 68 342 47 365 366 AOI222_X1 $T=49070 48600 0 180 $X=47435 $Y=47085
X2465 87 264 67 263 41 43 68 297 193 365 367 AOI222_X1 $T=50780 48600 0 0 $X=50665 $Y=48485
X2466 87 52 67 265 41 43 68 343 185 224 367 AOI222_X1 $T=54200 51400 0 180 $X=52565 $Y=49885
X2467 87 266 67 264 41 43 68 329 186 365 366 AOI222_X1 $T=53250 48600 1 0 $X=53135 $Y=47085
X2468 87 265 67 266 41 43 68 328 298 365 367 AOI222_X1 $T=56290 48600 1 180 $X=54655 $Y=48485
X2469 87 51 67 52 41 43 68 363 195 365 367 AOI222_X1 $T=56290 48600 0 0 $X=56175 $Y=48485
X2470 128 154 67 59 60 61 68 157 130 223 368 AOI222_X1 $T=62940 43000 0 0 $X=62825 $Y=42885
X2514 175 146 34 68 67 364 366 DLH_X1 $T=31970 45800 0 0 $X=31855 $Y=45685
X2515 43 176 261 68 67 364 368 DLH_X1 $T=44130 45800 1 0 $X=44015 $Y=44285
X2516 43 153 48 68 67 365 367 DLH_X1 $T=47170 48600 0 0 $X=47055 $Y=48485
X2517 43 127 260 68 67 223 368 DLH_X1 $T=47740 43000 0 0 $X=47625 $Y=42885
X2518 43 177 264 68 67 364 366 DLH_X1 $T=50210 45800 0 0 $X=50095 $Y=45685
X2519 43 88 263 68 67 364 368 DLH_X1 $T=50780 45800 1 0 $X=50665 $Y=44285
X2520 43 178 49 68 67 224 367 DLH_X1 $T=50780 51400 1 0 $X=50665 $Y=49885
X2521 43 154 265 68 67 364 366 DLH_X1 $T=52110 45800 0 0 $X=51995 $Y=45685
X2522 43 155 266 68 67 364 368 DLH_X1 $T=52680 45800 1 0 $X=52565 $Y=44285
X2523 115 343 50 68 67 364 366 DLH_X1 $T=54390 45800 0 0 $X=54275 $Y=45685
X2524 43 179 51 68 67 364 368 DLH_X1 $T=56860 45800 1 0 $X=56745 $Y=44285
X2525 43 59 53 68 67 365 366 DLH_X1 $T=57430 48600 1 0 $X=57315 $Y=47085
X2526 43 180 52 68 67 224 367 DLH_X1 $T=58190 51400 1 0 $X=58075 $Y=49885
X2527 115 363 54 68 67 364 366 DLH_X1 $T=58570 45800 0 0 $X=58455 $Y=45685
X2528 115 328 55 68 67 364 368 DLH_X1 $T=58760 45800 1 0 $X=58645 $Y=44285
X2529 115 329 267 68 67 365 366 DLH_X1 $T=61230 48600 0 180 $X=59215 $Y=47085
X2530 115 159 56 68 67 365 367 DLH_X1 $T=60280 48600 0 0 $X=60165 $Y=48485
X2531 115 296 57 68 67 364 368 DLH_X1 $T=60660 45800 1 0 $X=60545 $Y=44285
X2532 115 297 62 68 67 365 366 DLH_X1 $T=64270 48600 1 0 $X=64155 $Y=47085
X2533 115 188 270 68 67 224 367 DLH_X1 $T=64270 51400 1 0 $X=64155 $Y=49885
X2534 115 342 63 68 67 364 368 DLH_X1 $T=64650 45800 1 0 $X=64535 $Y=44285
X2535 77 67 105 107 68 76 223 368 NOR3_X1 $T=20760 43000 0 0 $X=20645 $Y=42885
X2555 79 11 310 67 232 348 68 365 367 OAI211_X1 $T=14300 48600 1 180 $X=13235 $Y=48485
X2557 27 68 67 172 365 367 CLKBUF_X3 $T=25700 48600 0 0 $X=25585 $Y=48485
X2558 330 2 135 273 68 67 365 367 AOI21_X1 $T=2140 48600 0 0 $X=2025 $Y=48485
X2559 69 131 119 225 68 67 364 366 AOI21_X1 $T=3660 45800 0 0 $X=3545 $Y=45685
X2560 347 10 310 309 68 67 365 367 AOI21_X1 $T=13350 48600 1 180 $X=12475 $Y=48485
X2561 122 12 236 332 68 67 364 368 AOI21_X1 $T=15060 45800 1 0 $X=14945 $Y=44285
X2562 145 13 359 280 68 67 364 368 AOI21_X1 $T=17530 45800 0 180 $X=16655 $Y=44285
X2563 122 14 349 335 68 67 364 366 AOI21_X1 $T=18480 45800 1 180 $X=17605 $Y=45685
X2564 122 3 319 336 68 67 365 367 AOI21_X1 $T=18670 48600 1 180 $X=17795 $Y=48485
X2565 122 15 320 337 68 67 365 366 AOI21_X1 $T=18480 48600 1 0 $X=18365 $Y=47085
X2566 122 16 321 183 68 67 224 367 AOI21_X1 $T=18480 51400 1 0 $X=18365 $Y=49885
X2567 104 17 350 284 68 67 365 367 AOI21_X1 $T=20380 48600 0 0 $X=20265 $Y=48485
X2568 31 238 237 338 68 67 365 366 AOI21_X1 $T=26650 48600 1 0 $X=26535 $Y=47085
X2569 318 14 338 288 68 67 365 367 AOI21_X1 $T=28170 48600 0 0 $X=28055 $Y=48485
X2570 353 246 202 361 68 67 364 368 AOI21_X1 $T=33300 45800 0 180 $X=32425 $Y=44285
X2571 292 253 291 362 68 67 365 366 AOI21_X1 $T=38810 48600 0 180 $X=37935 $Y=47085
X2572 191 42 355 293 68 67 224 367 AOI21_X1 $T=42230 51400 0 180 $X=41355 $Y=49885
X2575 118 2 67 91 300 302 68 223 368 AOI22_X1 $T=1950 43000 1 180 $X=885 $Y=42885
X2576 344 1 67 92 358 303 68 365 366 AOI22_X1 $T=1000 48600 1 0 $X=885 $Y=47085
X2577 119 2 67 91 331 304 68 364 368 AOI22_X1 $T=3850 45800 1 0 $X=3735 $Y=44285
X2578 69 198 67 92 304 70 68 365 366 AOI22_X1 $T=3850 48600 1 0 $X=3735 $Y=47085
X2579 138 91 67 2 345 304 68 365 367 AOI22_X1 $T=3850 48600 0 0 $X=3735 $Y=48485
X2580 275 1 67 92 139 71 68 224 367 AOI22_X1 $T=3850 51400 1 0 $X=3735 $Y=49885
X2581 331 73 67 93 231 274 68 364 368 AOI22_X1 $T=4800 45800 1 0 $X=4685 $Y=44285
X2582 135 73 67 93 346 345 68 365 367 AOI22_X1 $T=4800 48600 0 0 $X=4685 $Y=48485
X2583 274 73 67 93 305 72 68 223 368 AOI22_X1 $T=4990 43000 0 0 $X=4875 $Y=42885
X2584 331 93 67 73 234 306 68 364 366 AOI22_X1 $T=6130 45800 0 0 $X=6015 $Y=45685
X2585 345 73 67 93 308 306 68 365 366 AOI22_X1 $T=6130 48600 1 0 $X=6015 $Y=47085
X2586 74 140 67 164 275 6 68 364 366 AOI22_X1 $T=7080 45800 0 0 $X=6965 $Y=45685
X2587 74 9 67 4 344 6 68 364 368 AOI22_X1 $T=7270 45800 1 0 $X=7155 $Y=44285
X2588 74 131 67 3 71 6 68 224 367 AOI22_X1 $T=8220 51400 0 180 $X=7155 $Y=49885
X2589 74 141 67 14 307 6 68 365 367 AOI22_X1 $T=8410 48600 1 180 $X=7345 $Y=48485
X2590 74 165 67 12 166 6 68 365 366 AOI22_X1 $T=8220 48600 1 0 $X=8105 $Y=47085
X2591 74 7 67 15 303 6 68 365 367 AOI22_X1 $T=8410 48600 0 0 $X=8295 $Y=48485
X2592 227 10 67 95 226 308 68 365 366 AOI22_X1 $T=9170 48600 1 0 $X=9055 $Y=47085
X2593 305 95 67 10 228 229 68 223 368 AOI22_X1 $T=9740 43000 0 0 $X=9625 $Y=42885
X2594 346 95 67 11 232 122 68 365 367 AOI22_X1 $T=10690 48600 0 0 $X=10575 $Y=48485
X2595 276 10 67 95 230 231 68 364 368 AOI22_X1 $T=12020 45800 1 0 $X=11905 $Y=44285
X2596 277 10 67 95 233 234 68 364 366 AOI22_X1 $T=12400 45800 0 0 $X=12285 $Y=45685
X2597 121 142 67 98 229 311 68 223 368 AOI22_X1 $T=13920 43000 0 0 $X=13805 $Y=42885
X2598 359 98 67 142 276 311 68 364 368 AOI22_X1 $T=14110 45800 1 0 $X=13995 $Y=44285
X2599 278 142 67 98 347 279 68 365 367 AOI22_X1 $T=14300 48600 0 0 $X=14185 $Y=48485
X2600 359 142 67 98 277 312 68 364 366 AOI22_X1 $T=14490 45800 0 0 $X=14375 $Y=45685
X2601 278 98 67 142 227 312 68 365 366 AOI22_X1 $T=14490 48600 1 0 $X=14375 $Y=47085
X2602 143 98 67 142 167 279 68 224 367 AOI22_X1 $T=15440 51400 0 180 $X=14375 $Y=49885
X2603 333 13 67 75 312 334 68 364 366 AOI22_X1 $T=16390 45800 1 180 $X=15325 $Y=45685
X2604 350 13 67 75 143 99 68 224 367 AOI22_X1 $T=16390 51400 0 180 $X=15325 $Y=49885
X2605 168 13 67 75 311 333 68 223 368 AOI22_X1 $T=16390 43000 0 0 $X=16275 $Y=42885
X2606 334 13 67 75 279 281 68 365 367 AOI22_X1 $T=16960 48600 0 0 $X=16845 $Y=48485
X2607 281 13 67 75 169 100 68 224 367 AOI22_X1 $T=17530 51400 1 0 $X=17415 $Y=49885
X2608 76 102 67 77 168 144 68 223 368 AOI22_X1 $T=19430 43000 1 180 $X=18365 $Y=42885
X2609 76 101 67 77 333 282 68 364 366 AOI22_X1 $T=18480 45800 0 0 $X=18365 $Y=45685
X2610 76 103 67 77 145 104 68 364 368 AOI22_X1 $T=19240 45800 1 0 $X=19125 $Y=44285
X2611 316 17 67 77 170 106 68 224 367 AOI22_X1 $T=19620 51400 1 0 $X=19505 $Y=49885
X2612 184 77 67 17 18 317 68 224 367 AOI22_X1 $T=21710 51400 1 0 $X=21595 $Y=49885
X2613 171 77 67 17 315 286 68 365 367 AOI22_X1 $T=23420 48600 1 180 $X=22355 $Y=48485
X2614 25 109 67 31 316 21 68 365 366 AOI22_X1 $T=23990 48600 1 0 $X=23875 $Y=47085
X2615 25 102 67 33 286 21 68 365 367 AOI22_X1 $T=25700 48600 1 180 $X=24635 $Y=48485
X2616 25 101 67 36 173 21 68 224 367 AOI22_X1 $T=27030 51400 1 0 $X=26915 $Y=49885
X2617 25 103 67 35 317 21 68 365 367 AOI22_X1 $T=27220 48600 0 0 $X=27105 $Y=48485
X2618 245 240 67 174 242 148 68 223 368 AOI22_X1 $T=29690 43000 0 0 $X=29575 $Y=42885
X2619 33 244 67 360 288 323 68 224 367 AOI22_X1 $T=30640 51400 1 0 $X=30525 $Y=49885
X2620 290 3 67 15 323 322 68 365 367 AOI22_X1 $T=31970 48600 1 180 $X=30905 $Y=48485
X2621 257 327 67 339 254 325 68 365 366 AOI22_X1 $T=40710 48600 1 0 $X=40595 $Y=47085
X2622 128 59 67 178 156 89 68 223 368 AOI22_X1 $T=56480 43000 1 180 $X=55415 $Y=42885
X2623 129 157 67 153 199 60 68 223 368 AOI22_X1 $T=57810 43000 0 0 $X=57695 $Y=42885
X2624 89 59 67 157 299 60 68 223 368 AOI22_X1 $T=61990 43000 0 0 $X=61875 $Y=42885
X2625 120 1 68 137 92 303 67 224 367 OAI22_X1 $T=2520 51400 1 0 $X=2405 $Y=49885
X2626 347 97 68 309 96 346 67 365 367 OAI22_X1 $T=12590 48600 1 180 $X=11525 $Y=48485
X2627 245 240 68 289 243 324 67 364 368 OAI22_X1 $T=32540 45800 0 180 $X=31475 $Y=44285
X2628 339 325 68 326 241 256 67 364 366 OAI22_X1 $T=36340 45800 0 0 $X=36225 $Y=45685
X2629 257 327 68 354 348 352 67 365 367 OAI22_X1 $T=39000 48600 1 180 $X=37935 $Y=48485
X2630 113 152 68 114 84 83 67 224 367 OAI22_X1 $T=39570 51400 1 0 $X=39455 $Y=49885
X2631 308 96 68 226 227 67 97 336 365 366 OAI221_X1 $T=10120 48600 1 0 $X=10005 $Y=47085
X2632 305 96 68 228 229 67 97 332 223 368 OAI221_X1 $T=10690 43000 0 0 $X=10575 $Y=42885
X2633 276 97 68 230 231 67 96 335 223 368 OAI221_X1 $T=11830 43000 0 0 $X=11715 $Y=42885
X2634 277 97 68 233 234 67 96 337 364 366 OAI221_X1 $T=13350 45800 0 0 $X=13235 $Y=45685
X2635 287 12 68 237 26 67 164 201 223 368 OAI221_X1 $T=26080 43000 1 180 $X=24825 $Y=42885
X2636 166 1 302 301 68 67 364 368 OAI21_X1 $T=1000 45800 1 0 $X=885 $Y=44285
X2637 344 1 118 136 68 67 223 368 OAI21_X1 $T=1950 43000 0 0 $X=1835 $Y=42885
X2638 330 2 306 272 68 67 365 366 OAI21_X1 $T=1950 48600 1 0 $X=1835 $Y=47085
X2639 350 13 278 313 68 67 365 367 OAI21_X1 $T=16200 48600 0 0 $X=16085 $Y=48485
X2640 282 77 281 235 68 67 365 367 OAI21_X1 $T=19620 48600 0 0 $X=19505 $Y=48485
X2641 316 17 314 283 68 67 365 366 OAI21_X1 $T=20380 48600 1 0 $X=20265 $Y=47085
X2642 144 77 334 285 68 67 364 366 OAI21_X1 $T=21520 45800 0 0 $X=21405 $Y=45685
X2643 79 12 243 236 68 67 364 368 OAI21_X1 $T=24180 45800 0 180 $X=23305 $Y=44285
X2644 79 14 245 349 68 67 364 366 OAI21_X1 $T=24180 45800 0 0 $X=24065 $Y=45685
X2645 79 3 339 319 68 67 365 366 OAI21_X1 $T=29690 48600 0 180 $X=28815 $Y=47085
X2646 79 15 241 320 68 67 365 366 OAI21_X1 $T=29880 48600 1 0 $X=29765 $Y=47085
X2647 79 16 257 321 68 67 224 367 OAI21_X1 $T=29880 51400 1 0 $X=29765 $Y=49885
X2648 150 242 361 149 68 67 223 368 OAI21_X1 $T=31400 43000 1 180 $X=30525 $Y=42885
X2649 326 254 362 340 68 67 364 366 OAI21_X1 $T=38430 45800 0 0 $X=38315 $Y=45685
X2650 114 134 293 294 68 67 224 367 OAI21_X1 $T=42230 51400 1 0 $X=42115 $Y=49885
X2651 302 68 2 272 67 364 368 NAND2_X1 $T=1760 45800 1 0 $X=1645 $Y=44285
X2652 69 68 190 301 67 364 368 NAND2_X1 $T=2900 45800 0 180 $X=2215 $Y=44285
X2653 314 68 13 313 67 365 366 NAND2_X1 $T=17720 48600 0 180 $X=17035 $Y=47085
X2654 76 68 146 283 67 364 366 NAND2_X1 $T=21520 45800 1 180 $X=20835 $Y=45685
X2655 173 68 77 235 67 224 367 NAND2_X1 $T=21710 51400 0 180 $X=21025 $Y=49885
X2656 286 68 77 285 67 365 366 NAND2_X1 $T=23040 48600 0 180 $X=22355 $Y=47085
X2657 111 68 81 112 67 365 366 NAND2_X1 $T=35580 48600 1 0 $X=35465 $Y=47085
X2658 256 68 241 340 67 364 366 NAND2_X1 $T=39760 45800 1 180 $X=39075 $Y=45685
X2659 83 68 84 294 67 224 367 NAND2_X1 $T=44130 51400 0 180 $X=43445 $Y=49885
X2660 158 68 299 267 67 223 368 NAND2_X1 $T=60280 43000 0 0 $X=60165 $Y=42885
X2661 189 67 2 273 68 224 367 NOR2_X1 $T=1950 51400 1 0 $X=1835 $Y=49885
X2662 275 67 1 225 68 364 366 NOR2_X1 $T=4990 45800 1 180 $X=4305 $Y=45685
X2663 314 67 13 280 68 364 366 NOR2_X1 $T=17720 45800 1 180 $X=17035 $Y=45685
X2664 317 67 17 284 68 365 367 NOR2_X1 $T=22470 48600 1 180 $X=21785 $Y=48485
X2665 105 67 107 21 68 223 368 NOR2_X1 $T=22850 43000 0 0 $X=22735 $Y=42885
X2666 105 67 108 25 68 364 368 NOR2_X1 $T=23420 45800 0 180 $X=22735 $Y=44285
X2667 289 67 150 246 68 223 368 NOR2_X1 $T=31970 43000 1 180 $X=31285 $Y=42885
X2668 354 67 326 253 68 365 366 NOR2_X1 $T=38050 48600 0 180 $X=37365 $Y=47085
X2685 68 256 258 255 67 364 368 XNOR2_X1 $T=39190 45800 1 0 $X=39075 $Y=44285
X2686 68 241 260 258 67 223 368 XNOR2_X1 $T=39760 43000 0 0 $X=39645 $Y=42885
X2687 68 83 262 295 67 224 367 XNOR2_X1 $T=44130 51400 1 0 $X=44015 $Y=49885
X2688 68 84 266 262 67 365 367 XNOR2_X1 $T=47170 48600 1 180 $X=45915 $Y=48485
X2689 151 250 324 243 67 68 40 223 368 FA_X1 $T=35010 43000 1 180 $X=31855 $Y=42885
X2690 250 245 240 353 67 68 44 364 368 FA_X1 $T=33300 45800 1 0 $X=33185 $Y=44285
X2691 259 257 327 292 67 68 264 365 367 FA_X1 $T=39000 48600 0 0 $X=38885 $Y=48485
X2692 255 341 325 339 67 68 261 364 366 FA_X1 $T=39760 45800 0 0 $X=39645 $Y=45685
X2693 341 259 352 348 67 68 263 365 366 FA_X1 $T=41660 48600 1 0 $X=41545 $Y=47085
X2694 295 46 152 113 67 68 265 224 367 FA_X1 $T=45270 51400 1 0 $X=45155 $Y=49885
X2706 110 287 68 78 28 30 67 239 324 364 368 OAI222_X1 $T=26270 45800 1 0 $X=26155 $Y=44285
X2707 110 318 68 31 28 30 67 238 240 365 366 OAI222_X1 $T=28930 48600 0 180 $X=27295 $Y=47085
X2708 110 322 68 33 28 30 67 244 256 364 366 OAI222_X1 $T=30450 45800 0 0 $X=30335 $Y=45685
X2709 110 290 68 35 28 30 67 247 325 365 366 OAI222_X1 $T=33110 48600 1 0 $X=32995 $Y=47085
X2710 110 251 68 36 28 30 67 248 352 365 367 OAI222_X1 $T=35200 48600 1 180 $X=33565 $Y=48485
X2711 110 252 68 38 28 30 67 39 327 224 367 OAI222_X1 $T=37670 51400 1 0 $X=37555 $Y=49885
X2713 36 248 67 249 35 68 247 351 224 367 AOI221_X1 $T=33870 51400 0 180 $X=32615 $Y=49885
X2714 251 11 67 37 252 68 16 249 224 367 AOI221_X1 $T=35010 51400 1 0 $X=34895 $Y=49885
X2715 123 29 78 68 239 124 67 223 368 AOI211_X1 $T=27030 43000 0 0 $X=26915 $Y=42885
X2717 112 82 68 67 365 366 INV_X2 $T=36150 48600 1 0 $X=36035 $Y=47085
X2718 147 105 108 68 107 105 287 282 67 364 368 OAI33_X1 $T=21520 45800 0 180 $X=20075 $Y=44285
X2720 200 6 94 68 67 223 368 NOR2_X2 $T=7460 43000 0 0 $X=7345 $Y=42885
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 9 A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 10 A2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_10
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 249 250
** N=418 EP=243 IP=5837 FDC=2078
M0 3 109 104 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=7075 $Y=42495 $D=1
M1 104 8 3 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7265 $Y=42495 $D=1
M2 3 9 104 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7455 $Y=42495 $D=1
M3 104 9 3 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7645 $Y=42495 $D=1
M4 3 8 104 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=7835 $Y=42495 $D=1
M5 104 109 3 249 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=8025 $Y=42495 $D=1
M6 104 40 323 413 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=33295 $Y=39695 $D=1
M7 55 323 104 413 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=33485 $Y=39695 $D=1
M8 104 323 55 413 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=33675 $Y=39695 $D=1
M9 409 109 105 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=7075 $Y=41690 $D=0
M10 410 8 409 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7265 $Y=41690 $D=0
M11 3 9 410 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7455 $Y=41690 $D=0
M12 411 9 3 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7645 $Y=41690 $D=0
M13 412 8 411 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=7835 $Y=41690 $D=0
M14 105 109 412 416 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=8025 $Y=41690 $D=0
M15 105 40 323 417 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=33295 $Y=38890 $D=0
M16 55 323 105 417 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=33485 $Y=38890 $D=0
M17 105 323 55 417 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=33675 $Y=38890 $D=0
X2233 135 1 104 105 107 414 250 AND2_X1 $T=1000 34600 1 0 $X=885 $Y=33085
X2234 5 7 104 105 108 415 418 AND2_X1 $T=6890 37400 1 0 $X=6775 $Y=35885
X2235 9 142 104 105 216 249 416 AND2_X1 $T=8220 43000 1 0 $X=8105 $Y=41485
X2236 5 18 104 105 144 415 417 AND2_X1 $T=13920 37400 0 0 $X=13805 $Y=37285
X2237 135 62 104 105 284 414 418 AND2_X1 $T=45840 34600 0 0 $X=45725 $Y=34485
X2238 135 71 104 105 285 413 417 AND2_X1 $T=50780 40200 1 0 $X=50665 $Y=38685
X2239 75 292 104 105 304 413 417 AND2_X1 $T=52300 40200 0 180 $X=51425 $Y=38685
X2240 75 293 104 105 170 249 416 AND2_X1 $T=51920 43000 1 0 $X=51805 $Y=41485
X2241 135 190 104 105 221 249 416 AND2_X1 $T=52680 43000 1 0 $X=52565 $Y=41485
X2251 284 58 104 105 280 415 418 DFF_X1 $T=40900 37400 1 0 $X=40785 $Y=35885
X2252 285 58 104 105 281 413 416 DFF_X1 $T=41850 40200 0 0 $X=41735 $Y=40085
X2253 304 102 104 105 178 249 416 DFF_X1 $T=66170 43000 1 0 $X=66055 $Y=41485
X2833 193 104 105 2 414 418 INV_X1 $T=1570 34600 0 0 $X=1455 $Y=34485
X2834 22 104 105 136 414 250 INV_X1 $T=3280 34600 1 0 $X=3165 $Y=33085
X2835 137 104 105 264 414 250 INV_X1 $T=4610 34600 1 0 $X=4495 $Y=33085
X2836 140 104 105 139 413 417 INV_X1 $T=8030 40200 0 180 $X=7535 $Y=38685
X2837 387 104 105 339 415 417 INV_X1 $T=8030 37400 0 0 $X=7915 $Y=37285
X2838 142 104 105 8 413 416 INV_X1 $T=8410 40200 1 180 $X=7915 $Y=40085
X2839 342 104 105 340 415 418 INV_X1 $T=8410 37400 1 0 $X=8295 $Y=35885
X2840 385 104 105 341 414 418 INV_X1 $T=8980 34600 0 0 $X=8865 $Y=34485
X2841 373 104 105 343 414 418 INV_X1 $T=10120 34600 0 0 $X=10005 $Y=34485
X2842 11 104 105 143 415 417 INV_X1 $T=10310 37400 0 0 $X=10195 $Y=37285
X2843 25 104 105 182 413 416 INV_X1 $T=12590 40200 0 0 $X=12475 $Y=40085
X2844 218 104 105 14 413 417 INV_X1 $T=14300 40200 0 180 $X=13805 $Y=38685
X2845 110 104 105 198 249 416 INV_X1 $T=15630 43000 0 180 $X=15135 $Y=41485
X2846 26 104 105 353 414 418 INV_X1 $T=19240 34600 1 180 $X=18745 $Y=34485
X2847 112 104 105 23 414 250 INV_X1 $T=20570 34600 0 180 $X=20075 $Y=33085
X2848 116 104 105 401 415 418 INV_X1 $T=20190 37400 1 0 $X=20075 $Y=35885
X2849 156 104 105 153 413 417 INV_X1 $T=22850 40200 0 180 $X=22355 $Y=38685
X2850 152 104 105 114 249 416 INV_X1 $T=23230 43000 0 180 $X=22735 $Y=41485
X2851 117 104 105 262 415 417 INV_X1 $T=23230 37400 0 0 $X=23115 $Y=37285
X2852 115 104 105 267 413 417 INV_X1 $T=23420 40200 1 0 $X=23305 $Y=38685
X2853 30 104 105 183 414 250 INV_X1 $T=23990 34600 1 0 $X=23875 $Y=33085
X2854 34 104 105 271 413 416 INV_X1 $T=25510 40200 1 180 $X=25015 $Y=40085
X2855 150 104 105 269 415 418 INV_X1 $T=25890 37400 0 180 $X=25395 $Y=35885
X2856 33 104 105 266 414 418 INV_X1 $T=26080 34600 1 180 $X=25585 $Y=34485
X2857 27 104 105 184 414 250 INV_X1 $T=26270 34600 1 0 $X=26155 $Y=33085
X2858 119 104 105 272 413 417 INV_X1 $T=27220 40200 0 180 $X=26725 $Y=38685
X2859 20 104 105 273 413 416 INV_X1 $T=28360 40200 1 180 $X=27865 $Y=40085
X2860 32 104 105 38 249 416 INV_X1 $T=28360 43000 0 180 $X=27865 $Y=41485
X2861 208 104 105 274 415 417 INV_X1 $T=32540 37400 1 180 $X=32045 $Y=37285
X2862 229 104 105 324 414 418 INV_X1 $T=37670 34600 0 0 $X=37555 $Y=34485
X2863 406 104 105 325 415 417 INV_X1 $T=41280 37400 0 0 $X=41165 $Y=37285
X2864 326 104 105 293 415 417 INV_X1 $T=42800 37400 0 0 $X=42685 $Y=37285
X2865 231 104 105 292 414 418 INV_X1 $T=42990 34600 0 0 $X=42875 $Y=34485
X2866 82 104 105 64 415 417 INV_X1 $T=44320 37400 0 0 $X=44205 $Y=37285
X2867 407 104 105 327 413 416 INV_X1 $T=45080 40200 0 0 $X=44965 $Y=40085
X2868 68 104 105 191 414 418 INV_X1 $T=46600 34600 0 0 $X=46485 $Y=34485
X2869 360 104 105 164 414 250 INV_X1 $T=47550 34600 1 0 $X=47435 $Y=33085
X2870 332 104 105 365 413 417 INV_X1 $T=55530 40200 0 180 $X=55035 $Y=38685
X2871 84 104 105 67 413 416 INV_X1 $T=56670 40200 0 0 $X=56555 $Y=40085
X2872 93 104 105 66 414 418 INV_X1 $T=60470 34600 0 0 $X=60355 $Y=34485
X2873 174 104 105 176 415 417 INV_X1 $T=62370 37400 0 0 $X=62255 $Y=37285
X2874 192 104 105 89 414 418 INV_X1 $T=62940 34600 1 180 $X=62445 $Y=34485
X2875 69 104 105 73 414 418 INV_X1 $T=62940 34600 0 0 $X=62825 $Y=34485
X2876 85 104 105 92 415 418 INV_X1 $T=64460 37400 1 0 $X=64345 $Y=35885
X2877 177 104 105 76 415 417 INV_X1 $T=65790 37400 0 0 $X=65675 $Y=37285
X2878 86 104 105 103 414 250 INV_X1 $T=68260 34600 1 0 $X=68145 $Y=33085
X2879 101 104 105 171 413 417 INV_X1 $T=68450 40200 1 0 $X=68335 $Y=38685
X2880 98 104 105 91 413 417 INV_X1 $T=68830 40200 1 0 $X=68715 $Y=38685
X2954 401 262 105 14 351 16 104 117 261 415 417 AOI222_X1 $T=20190 37400 0 0 $X=20075 $Y=37285
X2955 401 267 105 14 263 16 104 115 318 415 418 AOI222_X1 $T=20570 37400 1 0 $X=20455 $Y=35885
X2956 319 358 105 31 30 26 104 264 260 414 250 AOI222_X1 $T=23610 34600 0 180 $X=21975 $Y=33085
X2957 226 46 105 48 280 50 104 324 326 415 418 AOI222_X1 $T=37290 37400 1 0 $X=37175 $Y=35885
X2958 126 282 105 283 52 51 104 377 235 413 417 AOI222_X1 $T=38050 40200 1 0 $X=37935 $Y=38685
X2959 126 53 105 282 52 51 104 376 225 249 416 AOI222_X1 $T=40330 43000 0 180 $X=38695 $Y=41485
X2960 226 54 105 48 281 55 104 325 187 413 416 AOI222_X1 $T=40330 40200 0 0 $X=40215 $Y=40085
X2961 126 61 105 56 52 57 104 403 406 414 250 AOI222_X1 $T=41470 34600 1 0 $X=41355 $Y=33085
X2962 126 283 105 61 52 51 104 378 407 415 418 AOI222_X1 $T=44130 37400 1 0 $X=44015 $Y=35885
X2963 226 45 105 48 49 55 104 327 232 413 416 AOI222_X1 $T=48120 40200 1 180 $X=46485 $Y=40085
X2964 87 72 105 68 67 64 104 162 394 415 417 AOI222_X1 $T=50970 37400 1 180 $X=49335 $Y=37285
X2965 70 85 105 86 64 87 104 101 382 413 416 AOI222_X1 $T=58190 40200 0 0 $X=58075 $Y=40085
X2966 64 88 105 63 73 87 104 162 236 414 250 AOI222_X1 $T=58950 34600 1 0 $X=58835 $Y=33085
X2967 89 86 105 93 70 73 104 99 227 414 250 AOI222_X1 $T=62750 34600 1 0 $X=62635 $Y=33085
X2968 215 94 105 85 96 95 104 98 334 414 250 AOI222_X1 $T=64270 34600 1 0 $X=64155 $Y=33085
X2969 96 98 105 97 95 81 104 85 370 415 417 AOI222_X1 $T=65790 37400 1 180 $X=64155 $Y=37285
X2970 87 86 105 80 64 81 104 97 301 415 417 AOI222_X1 $T=67880 37400 1 180 $X=66245 $Y=37285
X2971 87 80 105 93 67 64 104 74 405 413 417 AOI222_X1 $T=66930 40200 1 0 $X=66815 $Y=38685
X2972 87 93 105 74 67 64 104 63 371 415 417 AOI222_X1 $T=67880 37400 0 0 $X=67765 $Y=37285
X3025 50 115 189 104 105 415 418 DLH_X1 $T=29500 37400 0 180 $X=27485 $Y=35885
X3026 50 33 41 104 105 415 418 DLH_X1 $T=29500 37400 1 0 $X=29385 $Y=35885
X3027 55 34 45 104 105 413 417 DLH_X1 $T=33870 40200 1 0 $X=33755 $Y=38685
X3028 50 150 46 104 105 414 418 DLH_X1 $T=34060 34600 0 0 $X=33945 $Y=34485
X3029 55 117 280 104 105 415 417 DLH_X1 $T=34440 37400 0 0 $X=34325 $Y=37285
X3030 55 12 281 104 105 413 416 DLH_X1 $T=38050 40200 1 180 $X=36035 $Y=40085
X3031 55 20 49 104 105 249 416 DLH_X1 $T=36910 43000 1 0 $X=36795 $Y=41485
X3032 51 209 282 104 105 415 417 DLH_X1 $T=39190 37400 1 180 $X=37175 $Y=37285
X3033 57 88 283 104 105 414 250 DLH_X1 $T=39570 34600 1 0 $X=39455 $Y=33085
X3034 51 162 53 104 105 413 417 DLH_X1 $T=39570 40200 1 0 $X=39455 $Y=38685
X3035 166 403 59 104 105 414 250 DLH_X1 $T=42990 34600 1 0 $X=42875 $Y=33085
X3036 51 68 60 104 105 413 417 DLH_X1 $T=43560 40200 1 0 $X=43445 $Y=38685
X3037 166 378 286 104 105 415 418 DLH_X1 $T=45650 37400 1 0 $X=45535 $Y=35885
X3038 166 377 287 104 105 415 417 DLH_X1 $T=49450 37400 1 180 $X=47435 $Y=37285
X3039 166 167 65 104 105 413 417 DLH_X1 $T=48880 40200 1 0 $X=48765 $Y=38685
X3040 166 376 290 104 105 249 416 DLH_X1 $T=50020 43000 1 0 $X=49905 $Y=41485
X3041 166 169 294 104 105 413 416 DLH_X1 $T=52110 40200 0 0 $X=51995 $Y=40085
X3042 45 105 54 46 41 125 104 415 418 NOR4_X1 $T=34630 37400 1 0 $X=34515 $Y=35885
X3043 49 105 281 280 189 359 104 415 417 NOR4_X1 $T=37290 37400 1 180 $X=36225 $Y=37285
X3044 289 104 210 395 361 287 105 415 418 NAND4_X1 $T=50590 37400 1 0 $X=50475 $Y=35885
X3045 331 104 396 211 362 286 105 415 418 NAND4_X1 $T=54010 37400 1 0 $X=53895 $Y=35885
X3046 366 104 397 365 364 290 105 413 417 NAND4_X1 $T=55150 40200 0 180 $X=54085 $Y=38685
X3047 379 104 300 370 405 224 105 413 416 NAND4_X1 $T=63700 40200 0 0 $X=63585 $Y=40085
X3048 196 105 8 9 104 335 413 416 NOR3_X1 $T=6700 40200 0 0 $X=6585 $Y=40085
X3049 154 105 153 152 104 317 413 417 NOR3_X1 $T=21520 40200 0 180 $X=20645 $Y=38685
X3050 296 105 168 171 104 328 414 418 NOR3_X1 $T=50210 34600 1 180 $X=49335 $Y=34485
X3051 131 105 130 171 104 297 414 250 NOR3_X1 $T=56100 34600 0 180 $X=55225 $Y=33085
X3052 131 105 172 91 104 333 414 250 NOR3_X1 $T=56100 34600 1 0 $X=55985 $Y=33085
X3071 116 12 344 105 408 277 104 415 417 OAI211_X1 $T=11830 37400 1 180 $X=10765 $Y=37285
X3072 263 25 355 105 318 157 104 414 418 OAI211_X1 $T=19240 34600 0 0 $X=19125 $Y=34485
X3073 351 25 356 105 261 392 104 415 417 OAI211_X1 $T=19240 37400 0 0 $X=19125 $Y=37285
X3074 69 66 394 105 288 363 104 415 418 OAI211_X1 $T=50590 37400 0 180 $X=49525 $Y=35885
X3075 82 76 213 105 83 222 104 249 416 OAI211_X1 $T=55340 43000 1 0 $X=55225 $Y=41485
X3076 82 191 367 105 381 332 104 415 417 OAI211_X1 $T=58000 37400 1 180 $X=56935 $Y=37285
X3077 84 76 398 105 382 223 104 249 416 OAI211_X1 $T=58000 43000 1 0 $X=57885 $Y=41485
X3078 192 76 334 105 302 294 104 414 418 OAI211_X1 $T=64080 34600 0 0 $X=63965 $Y=34485
X3079 69 103 371 105 305 380 104 414 418 OAI211_X1 $T=69400 34600 1 180 $X=68335 $Y=34485
X3086 40 104 105 50 415 417 CLKBUF_X3 $T=29500 37400 0 0 $X=29385 $Y=37285
X3087 43 104 105 161 415 418 CLKBUF_X3 $T=31400 37400 1 0 $X=31285 $Y=35885
X3088 44 104 105 58 413 416 CLKBUF_X3 $T=31400 40200 0 0 $X=31285 $Y=40085
X3089 47 104 105 102 413 417 CLKBUF_X3 $T=35770 40200 1 0 $X=35655 $Y=38685
X3090 383 2 312 336 104 105 413 416 AOI21_X1 $T=2900 40200 1 180 $X=2025 $Y=40085
X3091 181 11 180 179 104 105 414 250 AOI21_X1 $T=11450 34600 0 180 $X=10575 $Y=33085
X3092 347 14 344 346 104 105 415 417 AOI21_X1 $T=12590 37400 1 180 $X=11715 $Y=37285
X3093 111 19 404 15 104 105 414 250 AOI21_X1 $T=14870 34600 1 0 $X=14755 $Y=33085
X3094 16 20 374 375 104 105 413 416 AOI21_X1 $T=15060 40200 0 0 $X=14945 $Y=40085
X3095 16 21 149 345 104 105 414 250 AOI21_X1 $T=17150 34600 1 0 $X=17035 $Y=33085
X3096 33 267 270 402 104 105 413 417 AOI21_X1 $T=25320 40200 1 0 $X=25205 $Y=38685
X3097 272 12 402 320 104 105 413 417 AOI21_X1 $T=26840 40200 0 180 $X=25965 $Y=38685
X3098 274 39 121 185 104 105 414 250 AOI21_X1 $T=29500 34600 0 180 $X=28625 $Y=33085
X3099 188 63 360 64 104 105 414 250 AOI21_X1 $T=46790 34600 1 0 $X=46675 $Y=33085
X3100 70 63 288 328 104 105 414 418 AOI21_X1 $T=48690 34600 0 0 $X=48575 $Y=34485
X3101 81 99 289 333 104 105 415 418 AOI21_X1 $T=54960 37400 1 0 $X=54845 $Y=35885
X3102 81 101 302 380 104 105 415 418 AOI21_X1 $T=65980 37400 1 0 $X=65865 $Y=35885
X3108 306 2 105 193 384 383 104 415 417 AOI22_X1 $T=1000 37400 0 0 $X=885 $Y=37285
X3109 3 22 105 117 383 335 104 413 417 AOI22_X1 $T=1000 40200 1 0 $X=885 $Y=38685
X3110 3 195 105 115 307 335 104 415 417 AOI22_X1 $T=3850 37400 1 180 $X=2785 $Y=37285
X3111 3 137 105 12 308 335 104 413 416 AOI22_X1 $T=3850 40200 1 180 $X=2785 $Y=40085
X3112 193 137 105 195 310 2 104 414 250 AOI22_X1 $T=4610 34600 0 180 $X=3545 $Y=33085
X3113 307 2 105 193 311 308 104 413 417 AOI22_X1 $T=3660 40200 1 0 $X=3545 $Y=38685
X3114 335 21 105 145 306 3 104 415 417 AOI22_X1 $T=3850 37400 0 0 $X=3735 $Y=37285
X3115 372 139 105 309 342 108 104 415 418 AOI22_X1 $T=5370 37400 0 180 $X=4305 $Y=35885
X3116 372 108 105 139 387 384 104 415 417 AOI22_X1 $T=4800 37400 0 0 $X=4685 $Y=37285
X3117 312 108 105 139 13 4 104 249 416 AOI22_X1 $T=5560 43000 1 0 $X=5445 $Y=41485
X3118 312 139 105 108 253 311 104 413 416 AOI22_X1 $T=5750 40200 0 0 $X=5635 $Y=40085
X3119 193 22 105 145 10 2 104 414 250 AOI22_X1 $T=6510 34600 1 0 $X=6395 $Y=33085
X3120 311 139 105 108 338 384 104 413 417 AOI22_X1 $T=6700 40200 1 0 $X=6585 $Y=38685
X3121 339 11 105 141 356 387 104 415 417 AOI22_X1 $T=8410 37400 0 0 $X=8295 $Y=37285
X3122 253 141 105 14 252 251 104 413 416 AOI22_X1 $T=9360 40200 1 180 $X=8295 $Y=40085
X3123 340 11 105 141 355 342 104 415 418 AOI22_X1 $T=8790 37400 1 0 $X=8675 $Y=35885
X3124 338 141 105 12 408 16 104 415 417 AOI22_X1 $T=9360 37400 0 0 $X=9245 $Y=37285
X3125 373 25 105 218 238 343 104 414 250 AOI22_X1 $T=9740 34600 1 0 $X=9625 $Y=33085
X3126 256 14 105 11 254 341 104 415 418 AOI22_X1 $T=11640 37400 0 180 $X=10575 $Y=35885
X3127 314 198 105 144 251 388 104 413 416 AOI22_X1 $T=12970 40200 0 0 $X=12855 $Y=40085
X3128 200 198 105 144 313 314 104 249 416 AOI22_X1 $T=13540 43000 1 0 $X=13425 $Y=41485
X3129 388 198 105 144 347 349 104 413 417 AOI22_X1 $T=14300 40200 1 0 $X=14185 $Y=38685
X3130 144 350 105 198 351 349 104 413 417 AOI22_X1 $T=15250 40200 1 0 $X=15135 $Y=38685
X3131 352 24 105 111 314 146 104 249 416 AOI22_X1 $T=15630 43000 1 0 $X=15515 $Y=41485
X3132 144 354 105 198 263 350 104 415 417 AOI22_X1 $T=16770 37400 1 180 $X=15705 $Y=37285
X3133 316 24 105 111 388 389 104 413 416 AOI22_X1 $T=15820 40200 0 0 $X=15705 $Y=40085
X3134 24 19 105 26 259 111 104 414 418 AOI22_X1 $T=16010 34600 0 0 $X=15895 $Y=34485
X3135 390 24 105 111 349 352 104 413 417 AOI22_X1 $T=17150 40200 0 180 $X=16085 $Y=38685
X3136 389 24 105 111 200 148 104 249 416 AOI22_X1 $T=16580 43000 1 0 $X=16465 $Y=41485
X3137 220 147 105 30 390 317 104 413 417 AOI22_X1 $T=19810 40200 0 180 $X=18745 $Y=38685
X3138 220 112 105 150 352 317 104 413 416 AOI22_X1 $T=19810 40200 1 180 $X=18745 $Y=40085
X3139 220 19 105 33 316 317 104 413 417 AOI22_X1 $T=19810 40200 1 0 $X=19695 $Y=38685
X3140 220 26 105 119 389 317 104 249 416 AOI22_X1 $T=19810 43000 1 0 $X=19695 $Y=41485
X3141 391 204 105 273 320 34 104 413 416 AOI22_X1 $T=25510 40200 0 0 $X=25395 $Y=40085
X3142 277 393 105 157 239 118 104 414 418 AOI22_X1 $T=28170 34600 1 180 $X=27105 $Y=34485
X3143 184 272 105 12 321 205 104 415 417 AOI22_X1 $T=28170 37400 1 180 $X=27105 $Y=37285
X3144 329 209 105 93 396 89 104 415 417 AOI22_X1 $T=53630 37400 0 0 $X=53515 $Y=37285
X3145 87 98 105 97 298 70 104 249 416 AOI22_X1 $T=54390 43000 1 0 $X=54275 $Y=41485
X3146 70 74 105 72 367 67 104 413 417 AOI22_X1 $T=57620 40200 0 180 $X=56555 $Y=38685
X3147 78 72 105 68 132 70 104 414 418 AOI22_X1 $T=56860 34600 0 0 $X=56745 $Y=34485
X3148 78 98 105 97 398 73 104 249 416 AOI22_X1 $T=59900 43000 0 180 $X=58835 $Y=41485
X3149 96 177 105 86 381 81 104 415 417 AOI22_X1 $T=60850 37400 1 180 $X=59785 $Y=37285
X3150 96 86 105 80 395 89 104 415 418 AOI22_X1 $T=60660 37400 1 0 $X=60545 $Y=35885
X3151 368 63 105 101 366 95 104 415 418 AOI22_X1 $T=61610 37400 1 0 $X=61495 $Y=35885
X3152 67 98 105 97 399 87 104 249 416 AOI22_X1 $T=62560 43000 0 180 $X=61495 $Y=41485
X3153 89 101 105 177 379 73 104 413 416 AOI22_X1 $T=62750 40200 0 0 $X=62635 $Y=40085
X3154 78 86 105 99 300 70 104 413 417 AOI22_X1 $T=63130 40200 1 0 $X=63015 $Y=38685
X3155 70 177 105 98 400 89 104 413 416 AOI22_X1 $T=64650 40200 0 0 $X=64535 $Y=40085
X3156 78 99 105 80 305 70 104 414 418 AOI22_X1 $T=67500 34600 0 0 $X=67385 $Y=34485
X3157 337 264 104 372 2 307 105 415 418 OAI22_X1 $T=2330 37400 1 0 $X=2215 $Y=35885
X3158 308 193 104 4 2 138 105 249 416 OAI22_X1 $T=3470 43000 1 0 $X=3355 $Y=41485
X3159 337 136 104 309 2 306 105 414 418 OAI22_X1 $T=3660 34600 0 0 $X=3545 $Y=34485
X3160 347 25 104 346 143 338 105 413 417 OAI22_X1 $T=12590 40200 0 180 $X=11525 $Y=38685
X3161 111 147 104 257 112 24 105 414 418 OAI22_X1 $T=16960 34600 0 0 $X=16845 $Y=34485
X3162 390 24 104 354 23 315 105 415 417 OAI22_X1 $T=18670 37400 1 180 $X=17605 $Y=37285
X3163 315 353 104 350 24 316 105 415 418 OAI22_X1 $T=17910 37400 1 0 $X=17795 $Y=35885
X3164 277 393 104 120 392 357 105 414 418 OAI22_X1 $T=28170 34600 0 0 $X=28055 $Y=34485
X3165 122 158 104 123 275 278 105 249 416 OAI22_X1 $T=29880 43000 1 0 $X=29765 $Y=41485
X3166 251 25 104 252 253 105 143 375 413 416 OAI221_X1 $T=9360 40200 0 0 $X=9245 $Y=40085
X3167 341 197 104 254 256 105 25 345 414 418 OAI221_X1 $T=11260 34600 0 0 $X=11145 $Y=34485
X3168 313 25 104 255 13 105 143 258 249 416 OAI221_X1 $T=11260 43000 1 0 $X=11145 $Y=41485
X3169 272 12 104 270 269 105 117 358 415 417 OAI221_X1 $T=25510 37400 1 180 $X=24255 $Y=37285
X3170 84 92 104 298 82 105 171 212 413 416 OAI221_X1 $T=56670 40200 1 180 $X=55415 $Y=40085
X3171 69 171 104 303 192 105 92 237 414 418 OAI221_X1 $T=66170 34600 1 180 $X=64915 $Y=34485
X3172 309 5 385 386 104 105 414 418 OAI21_X1 $T=5750 34600 0 0 $X=5635 $Y=34485
X3173 310 6 386 140 104 105 414 418 OAI21_X1 $T=6510 34600 0 0 $X=6395 $Y=34485
X3174 354 5 256 348 104 105 415 418 OAI21_X1 $T=12780 37400 1 0 $X=12665 $Y=35885
X3175 259 17 348 110 104 105 415 418 OAI21_X1 $T=13540 37400 1 0 $X=13425 $Y=35885
X3176 116 32 122 265 104 105 249 416 OAI21_X1 $T=23990 43000 0 180 $X=23115 $Y=41485
X3177 116 20 275 374 104 105 413 416 OAI21_X1 $T=24370 40200 0 0 $X=24255 $Y=40085
X3178 151 272 393 321 104 105 415 418 OAI21_X1 $T=26840 37400 1 0 $X=26725 $Y=35885
X3179 129 77 329 82 104 105 415 418 OAI21_X1 $T=53250 37400 1 0 $X=53135 $Y=35885
X3180 175 90 368 173 104 105 414 250 OAI21_X1 $T=61230 34600 0 180 $X=60355 $Y=33085
X3181 174 91 133 369 104 105 413 417 OAI21_X1 $T=60470 40200 1 0 $X=60355 $Y=38685
X3182 174 92 214 399 104 105 413 416 OAI21_X1 $T=61990 40200 0 0 $X=61875 $Y=40085
X3183 2 104 335 337 105 415 418 NAND2_X1 $T=1760 37400 1 0 $X=1645 $Y=35885
X3184 3 104 21 194 105 249 416 NAND2_X1 $T=3470 43000 0 180 $X=2785 $Y=41485
X3185 335 104 7 6 105 414 418 NAND2_X1 $T=7270 34600 0 0 $X=7155 $Y=34485
X3186 7 104 15 140 105 414 418 NAND2_X1 $T=8410 34600 1 180 $X=7725 $Y=34485
X3187 313 104 14 255 105 249 416 NAND2_X1 $T=11260 43000 0 180 $X=10575 $Y=41485
X3188 18 104 317 17 105 415 418 NAND2_X1 $T=14870 37400 1 0 $X=14755 $Y=35885
X3189 18 104 15 110 105 414 418 NAND2_X1 $T=16010 34600 1 180 $X=15325 $Y=34485
X3190 228 104 205 25 105 249 416 NAND2_X1 $T=17530 43000 1 0 $X=17415 $Y=41485
X3191 24 104 317 315 105 415 417 NAND2_X1 $T=18670 37400 0 0 $X=18555 $Y=37285
X3192 278 104 275 124 105 249 416 NAND2_X1 $T=30830 43000 1 0 $X=30715 $Y=41485
X3193 27 104 29 151 105 414 250 NAND2_X1 $T=34060 34600 1 0 $X=33945 $Y=33085
X3194 163 104 127 296 105 414 250 NAND2_X1 $T=44890 34600 1 0 $X=44775 $Y=33085
X3195 163 104 165 90 105 414 250 NAND2_X1 $T=47930 34600 1 0 $X=47815 $Y=33085
X3196 89 104 99 397 105 413 416 NAND2_X1 $T=54580 40200 1 180 $X=53895 $Y=40085
X3197 67 104 97 369 105 413 417 NAND2_X1 $T=61800 40200 0 180 $X=61115 $Y=38685
X3198 106 105 2 336 104 413 416 NOR2_X1 $T=1570 40200 0 0 $X=1455 $Y=40085
X3199 142 105 9 217 104 249 416 NOR2_X1 $T=8980 43000 1 0 $X=8865 $Y=41485
X3200 156 105 152 203 104 413 417 NOR2_X1 $T=22850 40200 1 0 $X=22735 $Y=38685
X3201 160 105 226 40 104 413 417 NOR2_X1 $T=30070 40200 0 180 $X=29385 $Y=38685
X3223 104 278 279 276 105 413 417 XNOR2_X1 $T=30830 40200 1 0 $X=30715 $Y=38685
X3224 104 275 283 279 105 413 417 XNOR2_X1 $T=33110 40200 0 180 $X=31855 $Y=38685
X3225 276 42 158 122 105 104 282 413 416 FA_X1 $T=31400 40200 1 180 $X=28245 $Y=40085
X3226 322 277 393 274 105 104 61 414 418 FA_X1 $T=32160 34600 1 180 $X=29005 $Y=34485
X3227 186 322 357 392 105 104 56 414 250 FA_X1 $T=32540 34600 0 180 $X=29385 $Y=33085
X3237 151 353 104 26 27 29 105 264 28 414 250 OAI222_X1 $T=20570 34600 1 0 $X=20455 $Y=33085
X3238 151 269 104 150 27 29 105 262 357 415 418 OAI222_X1 $T=25510 37400 0 180 $X=23875 $Y=35885
X3239 151 266 104 33 27 29 105 267 118 414 418 OAI222_X1 $T=24180 34600 0 0 $X=24065 $Y=34485
X3240 151 271 104 34 27 29 105 273 278 413 416 OAI222_X1 $T=26460 40200 0 0 $X=26345 $Y=40085
X3241 151 36 104 37 27 29 105 38 158 249 416 OAI222_X1 $T=26460 43000 1 0 $X=26345 $Y=41485
X3242 173 76 104 77 82 84 105 103 299 415 418 OAI222_X1 $T=56860 37400 1 0 $X=56745 $Y=35885
X3244 310 15 105 6 10 104 5 181 414 250 AOI221_X1 $T=7460 34600 1 0 $X=7345 $Y=33085
X3245 13 141 105 258 16 104 32 265 249 416 AOI221_X1 $T=12400 43000 1 0 $X=12285 $Y=41485
X3246 257 5 105 17 259 104 15 199 414 250 AOI221_X1 $T=12780 34600 1 0 $X=12665 $Y=33085
X3247 353 137 105 260 23 104 22 219 414 250 AOI221_X1 $T=19050 34600 0 180 $X=17795 $Y=33085
X3248 183 21 105 268 266 104 115 319 414 418 AOI221_X1 $T=24180 34600 1 180 $X=22925 $Y=34485
X3249 271 20 105 35 36 104 32 391 249 416 AOI221_X1 $T=25320 43000 1 0 $X=25205 $Y=41485
X3250 70 72 105 291 73 104 74 362 415 417 AOI221_X1 $T=50970 37400 0 0 $X=50855 $Y=37285
X3251 73 80 105 295 78 104 93 364 413 417 AOI221_X1 $T=53060 40200 1 0 $X=52945 $Y=38685
X3252 73 98 105 299 89 104 97 241 413 417 AOI221_X1 $T=59330 40200 1 0 $X=59215 $Y=38685
X3253 78 177 105 100 87 104 99 303 414 250 AOI221_X1 $T=66930 34600 0 180 $X=65675 $Y=33085
X3254 257 15 17 104 404 373 105 414 418 AOI211_X1 $T=12400 34600 0 0 $X=12285 $Y=34485
X3255 16 145 141 104 14 234 105 414 250 AOI211_X1 $T=16580 34600 0 180 $X=15515 $Y=33085
X3256 33 267 150 104 262 268 105 415 418 AOI211_X1 $T=23990 37400 0 180 $X=22925 $Y=35885
X3257 78 74 363 104 330 361 105 415 418 AOI211_X1 $T=51540 37400 1 0 $X=51425 $Y=35885
X3258 81 80 79 104 297 331 105 414 418 AOI211_X1 $T=54960 34600 1 180 $X=53895 $Y=34485
X3259 230 104 105 51 415 418 CLKBUF_X1 $T=39380 37400 0 180 $X=38695 $Y=35885
X3266 201 153 114 104 152 153 36 155 105 249 416 OAI33_X1 $T=22090 43000 0 180 $X=20645 $Y=41485
X3267 113 153 114 104 152 153 271 202 105 413 416 OAI33_X1 $T=22280 40200 0 0 $X=22165 $Y=40085
X3268 90 168 76 104 103 128 296 291 105 414 250 OAI33_X1 $T=50590 34600 1 0 $X=50475 $Y=33085
X3269 90 130 92 104 76 128 129 330 105 414 250 OAI33_X1 $T=51920 34600 1 0 $X=51805 $Y=33085
X3270 92 129 168 104 130 296 91 295 105 414 418 OAI33_X1 $T=52680 34600 0 0 $X=52565 $Y=34485
X3272 64 78 240 104 105 414 250 NOR2_X2 $T=48500 34600 1 0 $X=48385 $Y=33085
X3274 359 104 206 207 105 159 413 417 NAND3_X1 $T=28740 40200 1 0 $X=28625 $Y=38685
X3275 233 104 400 301 105 134 249 416 NAND3_X1 $T=64270 43000 1 0 $X=64155 $Y=41485
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 VSS VDD ZN 8 9
** N=13 EP=9 IP=0 FDC=10
M0 11 A1 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 12 A2 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 13 A3 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 10 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 10 A1 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD A2 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 10 A3 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 10 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X2 VSS A B VDD ZN 6 7
** N=12 EP=7 IP=0 FDC=16
M0 8 9 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=155 $Y=90 $D=1
M1 VSS 9 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=345 $Y=90 $D=1
M2 12 B VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=535 $Y=90 $D=1
M3 9 A 12 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=725 $Y=90 $D=1
M4 8 A ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=1110 $Y=90 $D=1
M5 ZN A 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1300 $Y=90 $D=1
M6 8 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=1490 $Y=90 $D=1
M7 ZN B 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1680 $Y=90 $D=1
M8 ZN 9 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=155 $Y=680 $D=0
M9 VDD 9 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=345 $Y=680 $D=0
M10 9 B VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=535 $Y=680 $D=0
M11 VDD A 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=725 $Y=680 $D=0
M12 ZN A 10 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=1110 $Y=680 $D=0
M13 11 A ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1300 $Y=680 $D=0
M14 VDD B 11 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=1490 $Y=680 $D=0
M15 10 B VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1680 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 262 263
** N=409 EP=239 IP=4808 FDC=1746
M0 403 26 96 405 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=15800 $Y=25695 $D=1
M1 31 21 403 405 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15990 $Y=25695 $D=1
M2 404 21 31 405 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16180 $Y=25695 $D=1
M3 96 26 404 405 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=16370 $Y=25695 $D=1
M4 96 331 332 406 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=48835 $Y=31890 $D=1
M5 332 292 96 406 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=49025 $Y=31890 $D=1
M6 96 62 332 406 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=49215 $Y=31890 $D=1
M7 284 332 96 406 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=49405 $Y=31890 $D=1
M8 31 26 95 262 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=15800 $Y=24890 $D=0
M9 95 21 31 262 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15990 $Y=24890 $D=0
M10 31 21 95 262 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16180 $Y=24890 $D=0
M11 95 26 31 262 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=16370 $Y=24890 $D=0
M12 401 331 332 263 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=48835 $Y=32795 $D=0
M13 402 292 401 263 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=49025 $Y=32795 $D=0
M14 95 62 402 263 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=49215 $Y=32795 $D=0
M15 284 332 95 263 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=49405 $Y=32480 $D=0
X1793 135 1 96 95 366 405 408 AND2_X1 $T=1000 26200 0 0 $X=885 $Y=26085
X1794 135 2 96 95 264 407 408 AND2_X1 $T=1760 29000 1 0 $X=1645 $Y=27485
X1795 136 5 96 95 343 405 262 AND2_X1 $T=5940 26200 1 0 $X=5825 $Y=24685
X1796 286 50 96 95 293 406 409 AND2_X1 $T=43560 31800 1 0 $X=43445 $Y=30285
X1797 358 50 96 95 55 406 263 AND2_X1 $T=43940 31800 0 0 $X=43825 $Y=31685
X1798 358 288 96 95 117 406 263 AND2_X1 $T=45650 31800 0 0 $X=45535 $Y=31685
X1799 92 86 96 95 340 405 262 AND2_X1 $T=64650 26200 0 180 $X=63775 $Y=24685
X1817 264 3 96 95 4 407 409 DFF_X1 $T=1000 29000 0 0 $X=885 $Y=28885
X1818 211 3 96 95 265 406 263 DFF_X1 $T=1000 31800 0 0 $X=885 $Y=31685
X1819 366 3 96 95 6 405 408 DFF_X1 $T=1760 26200 0 0 $X=1645 $Y=26085
X1820 343 8 96 95 24 405 262 DFF_X1 $T=6700 26200 1 0 $X=6585 $Y=24685
X2308 97 96 95 185 407 408 INV_X1 $T=9170 29000 1 0 $X=9055 $Y=27485
X2309 141 96 95 11 406 263 INV_X1 $T=9740 31800 0 0 $X=9625 $Y=31685
X2310 7 96 95 266 407 409 INV_X1 $T=14110 29000 0 0 $X=13995 $Y=28885
X2311 178 96 95 22 407 408 INV_X1 $T=16200 29000 1 0 $X=16085 $Y=27485
X2312 399 96 95 368 406 409 INV_X1 $T=18670 31800 0 180 $X=18175 $Y=30285
X2313 143 96 95 316 406 409 INV_X1 $T=18670 31800 1 0 $X=18555 $Y=30285
X2314 26 96 95 271 405 408 INV_X1 $T=19620 26200 0 0 $X=19505 $Y=26085
X2315 23 96 95 19 406 263 INV_X1 $T=19620 31800 0 0 $X=19505 $Y=31685
X2316 318 96 95 315 405 262 INV_X1 $T=20950 26200 1 0 $X=20835 $Y=24685
X2317 144 96 95 214 405 262 INV_X1 $T=21330 26200 1 0 $X=21215 $Y=24685
X2318 320 96 95 272 407 408 INV_X1 $T=22470 29000 0 180 $X=21975 $Y=27485
X2319 34 96 95 193 406 263 INV_X1 $T=23420 31800 0 0 $X=23305 $Y=31685
X2320 107 96 95 192 406 409 INV_X1 $T=23990 31800 1 0 $X=23875 $Y=30285
X2321 323 96 95 179 405 262 INV_X1 $T=27980 26200 1 0 $X=27865 $Y=24685
X2322 230 96 95 369 406 409 INV_X1 $T=29120 31800 0 180 $X=28625 $Y=30285
X2323 108 96 95 223 407 408 INV_X1 $T=31210 29000 1 0 $X=31095 $Y=27485
X2324 354 96 95 324 406 409 INV_X1 $T=35770 31800 1 0 $X=35655 $Y=30285
X2325 52 96 95 49 405 262 INV_X1 $T=38050 26200 1 0 $X=37935 $Y=24685
X2326 48 96 95 45 405 408 INV_X1 $T=38050 26200 0 0 $X=37935 $Y=26085
X2327 285 96 95 327 407 408 INV_X1 $T=41280 29000 0 180 $X=40785 $Y=27485
X2328 112 96 95 162 407 408 INV_X1 $T=41280 29000 1 0 $X=41165 $Y=27485
X2329 158 96 95 286 407 408 INV_X1 $T=41660 29000 1 0 $X=41545 $Y=27485
X2330 118 96 95 398 405 262 INV_X1 $T=48690 26200 1 0 $X=48575 $Y=24685
X2331 387 96 95 333 407 408 INV_X1 $T=50970 29000 0 180 $X=50475 $Y=27485
X2332 335 96 95 337 406 409 INV_X1 $T=53820 31800 1 0 $X=53705 $Y=30285
X2333 308 96 95 209 406 263 INV_X1 $T=63890 31800 0 0 $X=63775 $Y=31685
X2334 166 96 95 87 407 409 INV_X1 $T=65980 29000 1 180 $X=65485 $Y=28885
X2335 71 96 95 72 407 408 INV_X1 $T=66170 29000 1 0 $X=66055 $Y=27485
X2336 133 96 95 184 407 408 INV_X1 $T=68070 29000 1 0 $X=67955 $Y=27485
X2393 108 186 95 13 265 14 96 315 177 405 408 AOI222_X1 $T=11260 26200 0 0 $X=11145 $Y=26085
X2394 222 279 95 42 39 40 96 41 318 405 262 AOI222_X1 $T=29690 26200 1 0 $X=29575 $Y=24685
X2395 222 281 95 279 39 40 96 394 323 405 408 AOI222_X1 $T=31400 26200 0 0 $X=31285 $Y=26085
X2396 108 226 95 13 44 14 96 324 109 406 263 AOI222_X1 $T=34820 31800 0 0 $X=34705 $Y=31685
X2397 222 283 95 281 39 40 96 382 354 407 409 AOI222_X1 $T=35770 29000 0 0 $X=35655 $Y=28885
X2398 222 47 95 283 39 40 96 383 234 406 263 AOI222_X1 $T=38050 31800 0 0 $X=37935 $Y=31685
X2399 113 327 95 52 129 53 96 56 396 407 408 AOI222_X1 $T=44510 29000 1 0 $X=44395 $Y=27485
X2400 129 165 95 92 53 89 96 94 314 406 263 AOI222_X1 $T=69400 31800 1 180 $X=67765 $Y=31685
X2452 14 15 4 96 95 407 409 DLH_X1 $T=4230 29000 0 0 $X=4115 $Y=28885
X2453 14 16 265 96 95 406 409 DLH_X1 $T=4420 31800 1 0 $X=4305 $Y=30285
X2454 14 34 6 96 95 407 409 DLH_X1 $T=6130 29000 0 0 $X=6015 $Y=28885
X2455 14 7 9 96 95 405 408 DLH_X1 $T=8410 26200 0 0 $X=8295 $Y=26085
X2456 14 23 17 96 95 407 408 DLH_X1 $T=12970 29000 1 0 $X=12855 $Y=27485
X2457 14 213 186 96 95 405 408 DLH_X1 $T=18670 26200 1 180 $X=16655 $Y=26085
X2458 14 28 24 96 95 405 262 DLH_X1 $T=17720 26200 1 0 $X=17605 $Y=24685
X2459 14 35 30 96 95 405 408 DLH_X1 $T=20000 26200 0 0 $X=19885 $Y=26085
X2460 40 116 42 96 95 405 262 DLH_X1 $T=31210 26200 1 0 $X=31095 $Y=24685
X2461 40 180 279 96 95 407 408 DLH_X1 $T=31590 29000 1 0 $X=31475 $Y=27485
X2462 40 154 281 96 95 407 408 DLH_X1 $T=35390 29000 0 180 $X=33375 $Y=27485
X2463 156 394 373 96 95 405 262 DLH_X1 $T=36150 26200 1 0 $X=36035 $Y=24685
X2464 156 382 282 96 95 407 408 DLH_X1 $T=36340 29000 1 0 $X=36225 $Y=27485
X2465 40 52 283 96 95 407 409 DLH_X1 $T=37290 29000 0 0 $X=37175 $Y=28885
X2466 40 48 47 96 95 407 409 DLH_X1 $T=39190 29000 0 0 $X=39075 $Y=28885
X2467 156 383 284 96 95 406 263 DLH_X1 $T=39570 31800 0 0 $X=39455 $Y=31685
X2468 40 64 187 96 95 406 263 DLH_X1 $T=43370 31800 1 180 $X=41355 $Y=31685
X2469 6 95 265 4 9 375 96 405 408 NOR4_X1 $T=11260 26200 1 180 $X=10195 $Y=26085
X2470 115 95 51 291 180 328 96 407 409 NOR4_X1 $T=45270 29000 0 0 $X=45155 $Y=28885
X2471 202 95 361 385 301 360 96 405 408 NOR4_X1 $T=53820 26200 0 0 $X=53705 $Y=26085
X2472 123 95 90 235 125 361 96 405 262 NOR4_X1 $T=54200 26200 1 0 $X=54085 $Y=24685
X2473 120 95 90 81 171 390 96 407 408 NOR4_X1 $T=61040 29000 1 0 $X=60925 $Y=27485
X2474 201 96 128 293 162 217 95 407 409 NAND4_X1 $T=50210 29000 1 180 $X=49145 $Y=28885
X2475 388 96 337 203 300 68 95 406 263 NAND4_X1 $T=55340 31800 1 180 $X=54275 $Y=31685
X2476 128 96 170 88 72 400 95 407 409 NAND4_X1 $T=65980 29000 0 0 $X=65865 $Y=28885
X2477 112 95 158 57 96 325 405 408 NOR3_X1 $T=42420 26200 0 0 $X=42305 $Y=26085
X2478 326 95 66 88 96 386 406 263 NOR3_X1 $T=52110 31800 1 180 $X=51235 $Y=31685
X2479 170 95 66 298 96 336 407 409 NOR3_X1 $T=53630 29000 0 0 $X=53515 $Y=28885
X2480 362 95 336 302 96 300 407 409 NOR3_X1 $T=55150 29000 1 180 $X=54275 $Y=28885
X2481 88 95 169 133 96 303 406 409 NOR3_X1 $T=56480 31800 1 0 $X=56365 $Y=30285
X2482 118 95 77 81 96 304 407 408 NOR3_X1 $T=60090 29000 0 180 $X=59215 $Y=27485
X2498 100 7 376 95 268 145 96 407 408 OAI211_X1 $T=12970 29000 0 180 $X=11905 $Y=27485
X2499 100 16 139 95 270 278 96 406 263 OAI211_X1 $T=12780 31800 0 0 $X=12665 $Y=31685
X2500 391 75 76 95 79 389 96 406 263 OAI211_X1 $T=58950 31800 0 0 $X=58835 $Y=31685
X2501 74 78 363 95 307 305 96 406 409 OAI211_X1 $T=59330 31800 1 0 $X=59215 $Y=30285
X2502 74 84 364 95 85 208 96 406 263 OAI211_X1 $T=61420 31800 0 0 $X=61305 $Y=31685
X2505 138 7 397 185 96 95 406 409 AOI21_X1 $T=8030 31800 0 180 $X=7155 $Y=30285
X2506 344 10 267 220 96 95 406 409 AOI21_X1 $T=9360 31800 1 0 $X=9245 $Y=30285
X2507 212 269 268 346 96 95 406 409 AOI21_X1 $T=12590 31800 0 180 $X=11715 $Y=30285
X2508 101 15 367 393 96 95 407 409 AOI21_X1 $T=12590 29000 0 0 $X=12475 $Y=28885
X2509 369 274 320 321 96 95 407 409 AOI21_X1 $T=23610 29000 0 0 $X=23495 $Y=28885
X2510 287 46 357 180 96 95 407 408 AOI21_X1 $T=38810 29000 1 0 $X=38695 $Y=27485
X2511 398 51 224 325 96 95 405 262 AOI21_X1 $T=44510 26200 0 180 $X=43635 $Y=24685
X2512 58 54 290 45 96 95 407 408 AOI21_X1 $T=46030 29000 1 0 $X=45915 $Y=27485
X2513 119 291 331 69 96 95 406 409 AOI21_X1 $T=48880 31800 0 180 $X=48005 $Y=30285
X2514 124 299 335 80 96 95 407 408 AOI21_X1 $T=53820 29000 1 0 $X=53705 $Y=27485
X2515 123 58 302 69 96 95 407 408 AOI21_X1 $T=54580 29000 1 0 $X=54465 $Y=27485
X2516 339 80 182 88 96 95 405 408 AOI21_X1 $T=59520 26200 0 0 $X=59405 $Y=26085
X2517 82 83 307 390 96 95 407 409 AOI21_X1 $T=61420 29000 0 0 $X=61305 $Y=28885
X2518 131 84 372 210 96 95 405 408 AOI21_X1 $T=65410 26200 0 0 $X=65295 $Y=26085
X2520 10 345 95 7 376 101 96 407 409 AOI22_X1 $T=10690 29000 0 0 $X=10575 $Y=28885
X2521 189 212 95 16 270 101 96 406 263 AOI22_X1 $T=13730 31800 0 0 $X=13615 $Y=31685
X2522 19 7 95 107 317 22 96 406 409 AOI22_X1 $T=16010 31800 1 0 $X=15895 $Y=30285
X2523 178 192 95 368 378 317 96 407 409 AOI22_X1 $T=16770 29000 0 0 $X=16655 $Y=28885
X2524 278 104 95 145 276 105 96 407 409 AOI22_X1 $T=21520 29000 0 0 $X=21405 $Y=28885
X2525 216 70 95 161 215 356 96 405 262 AOI22_X1 $T=46980 26200 0 180 $X=45915 $Y=24685
X2526 129 83 95 70 313 89 96 407 408 AOI22_X1 $T=63510 29000 1 0 $X=63395 $Y=27485
X2527 189 140 96 190 11 98 95 406 263 OAI22_X1 $T=10120 31800 0 0 $X=10005 $Y=31685
X2528 269 140 96 346 11 345 95 406 409 OAI22_X1 $T=11830 31800 0 180 $X=10765 $Y=30285
X2529 145 105 96 350 148 106 95 405 408 OAI22_X1 $T=23420 26200 0 0 $X=23305 $Y=26085
X2530 278 104 96 275 377 322 95 407 409 OAI22_X1 $T=26460 29000 1 180 $X=25395 $Y=28885
X2531 149 153 96 353 349 379 95 406 409 OAI22_X1 $T=26650 31800 1 0 $X=26535 $Y=30285
X2532 58 157 96 338 78 119 95 405 408 OAI22_X1 $T=57810 26200 0 0 $X=57695 $Y=26085
X2533 29 192 96 31 36 95 107 106 406 409 OAI221_X1 $T=24370 31800 1 0 $X=24255 $Y=30285
X2534 121 65 96 295 294 95 120 373 405 262 OAI221_X1 $T=52110 26200 0 180 $X=50855 $Y=24685
X2535 119 72 96 313 87 95 170 311 407 409 OAI221_X1 $T=64460 29000 0 0 $X=64345 $Y=28885
X2536 308 69 96 314 87 95 204 219 406 409 OAI221_X1 $T=66740 31800 1 0 $X=66625 $Y=30285
X2538 344 11 393 267 96 95 406 409 OAI21_X1 $T=10120 31800 1 0 $X=10005 $Y=30285
X2539 22 12 347 138 96 95 407 408 OAI21_X1 $T=11260 29000 1 0 $X=11145 $Y=27485
X2540 100 15 377 367 96 95 407 409 OAI21_X1 $T=15250 29000 1 180 $X=14375 $Y=28885
X2541 192 20 348 99 96 95 407 409 OAI21_X1 $T=16770 29000 1 180 $X=15895 $Y=28885
X2542 100 22 148 142 96 95 407 408 OAI21_X1 $T=17340 29000 0 180 $X=16465 $Y=27485
X2543 271 272 103 143 96 95 407 408 OAI21_X1 $T=20950 29000 1 0 $X=20835 $Y=27485
X2544 100 34 349 146 96 95 406 409 OAI21_X1 $T=23230 31800 1 0 $X=23115 $Y=30285
X2545 350 276 321 351 96 95 407 408 OAI21_X1 $T=24560 29000 1 0 $X=24445 $Y=27485
X2546 353 37 221 352 96 95 406 263 OAI21_X1 $T=27980 31800 1 180 $X=27105 $Y=31685
X2547 357 45 356 355 96 95 405 262 OAI21_X1 $T=39190 26200 0 180 $X=38315 $Y=24685
X2548 328 289 198 83 96 95 407 409 OAI21_X1 $T=46220 29000 0 0 $X=46105 $Y=28885
X2549 298 60 330 200 96 95 407 409 OAI21_X1 $T=49260 29000 1 180 $X=48385 $Y=28885
X2550 163 60 164 119 96 95 405 262 OAI21_X1 $T=49070 26200 1 0 $X=48955 $Y=24685
X2551 163 72 371 58 96 95 407 408 OAI21_X1 $T=57240 29000 1 0 $X=57125 $Y=27485
X2552 171 60 374 341 96 95 405 408 OAI21_X1 $T=62750 26200 0 0 $X=62635 $Y=26085
X2553 372 88 183 342 96 95 405 262 OAI21_X1 $T=65790 26200 1 0 $X=65675 $Y=24685
X2554 90 92 392 170 96 95 405 408 OAI21_X1 $T=69400 26200 1 180 $X=68525 $Y=26085
X2555 316 96 229 140 95 406 409 NAND2_X1 $T=15440 31800 1 0 $X=15325 $Y=30285
X2556 319 96 271 100 95 407 409 NAND2_X1 $T=21140 29000 1 180 $X=20455 $Y=28885
X2557 106 96 148 351 95 407 408 NAND2_X1 $T=25890 29000 0 180 $X=25205 $Y=27485
X2558 379 96 349 352 95 406 263 NAND2_X1 $T=26650 31800 0 0 $X=26535 $Y=31685
X2559 45 96 49 285 95 405 408 NAND2_X1 $T=38430 26200 0 0 $X=38315 $Y=26085
X2560 384 96 155 355 95 405 262 NAND2_X1 $T=39760 26200 0 180 $X=39075 $Y=24685
X2561 56 96 57 110 95 405 262 NAND2_X1 $T=40900 26200 1 0 $X=40785 $Y=24685
X2562 358 96 286 181 95 407 408 NAND2_X1 $T=42040 29000 1 0 $X=41925 $Y=27485
X2563 293 96 287 326 95 407 409 NAND2_X1 $T=43940 29000 1 180 $X=43255 $Y=28885
X2564 327 96 293 169 95 407 409 NAND2_X1 $T=44510 29000 1 180 $X=43825 $Y=28885
X2565 293 96 358 120 95 406 409 NAND2_X1 $T=44320 31800 1 0 $X=44205 $Y=30285
X2566 114 96 116 58 95 405 408 NAND2_X1 $T=45270 26200 0 0 $X=45155 $Y=26085
X2567 288 96 55 199 95 406 263 NAND2_X1 $T=46410 31800 0 0 $X=46295 $Y=31685
X2568 288 96 52 200 95 407 409 NAND2_X1 $T=46980 29000 0 0 $X=46865 $Y=28885
X2569 293 96 162 298 95 406 409 NAND2_X1 $T=49450 31800 0 180 $X=48765 $Y=30285
X2570 359 96 370 292 95 406 409 NAND2_X1 $T=49450 31800 1 0 $X=49335 $Y=30285
X2571 122 96 94 123 95 405 408 NAND2_X1 $T=53250 26200 0 0 $X=53135 $Y=26085
X2572 88 96 93 218 95 405 262 NAND2_X1 $T=56860 26200 1 0 $X=56745 $Y=24685
X2573 53 96 115 363 95 406 263 NAND2_X1 $T=59900 31800 0 0 $X=59785 $Y=31685
X2574 127 96 128 77 95 405 408 NAND2_X1 $T=60850 26200 1 180 $X=60165 $Y=26085
X2575 122 96 128 308 95 407 409 NAND2_X1 $T=62750 29000 1 180 $X=62065 $Y=28885
X2576 233 96 130 341 95 405 408 NAND2_X1 $T=63510 26200 0 0 $X=63395 $Y=26085
X2577 132 96 210 391 95 405 408 NAND2_X1 $T=66740 26200 1 180 $X=66055 $Y=26085
X2578 316 95 21 10 96 406 409 NOR2_X1 $T=13920 31800 1 0 $X=13805 $Y=30285
X2579 143 95 378 319 96 407 408 NOR2_X1 $T=18670 29000 1 0 $X=18555 $Y=27485
X2580 275 95 350 274 96 407 408 NOR2_X1 $T=24560 29000 0 180 $X=23875 $Y=27485
X2581 196 95 353 194 96 406 263 NOR2_X1 $T=28550 31800 1 180 $X=27865 $Y=31685
X2582 39 95 231 43 96 405 408 NOR2_X1 $T=33490 26200 0 0 $X=33375 $Y=26085
X2583 52 95 154 287 96 407 408 NOR2_X1 $T=38240 29000 1 0 $X=38125 $Y=27485
X2584 112 95 52 358 96 407 409 NOR2_X1 $T=41090 29000 0 0 $X=40975 $Y=28885
X2585 56 95 64 50 96 406 263 NOR2_X1 $T=43940 31800 1 180 $X=43255 $Y=31685
X2586 160 95 116 288 96 405 262 NOR2_X1 $T=46030 26200 0 180 $X=45345 $Y=24685
X2587 326 95 69 289 96 406 409 NOR2_X1 $T=45650 31800 1 0 $X=45535 $Y=30285
X2588 299 95 129 166 96 405 408 NOR2_X1 $T=54770 26200 0 0 $X=54655 $Y=26085
X2589 120 95 69 172 96 407 408 NOR2_X1 $T=61990 29000 1 0 $X=61875 $Y=27485
X2590 199 95 66 312 96 406 263 NOR2_X1 $T=62370 31800 0 0 $X=62255 $Y=31685
X2591 91 95 120 173 96 406 409 NOR2_X1 $T=63320 31800 1 0 $X=63205 $Y=30285
X2613 96 379 280 277 95 406 409 XNOR2_X1 $T=27600 31800 1 0 $X=27485 $Y=30285
X2614 96 349 281 280 95 407 409 XNOR2_X1 $T=30640 29000 1 180 $X=29385 $Y=28885
X2615 33 273 322 377 95 96 42 405 262 FA_X1 $T=21710 26200 1 0 $X=21595 $Y=24685
X2616 273 278 104 369 95 96 279 407 409 FA_X1 $T=29500 29000 1 180 $X=26345 $Y=28885
X2617 277 38 153 149 95 96 283 406 409 FA_X1 $T=29120 31800 1 0 $X=29005 $Y=30285
X2622 102 27 96 28 29 31 95 32 322 406 263 OAI222_X1 $T=20000 31800 0 0 $X=19885 $Y=31685
X2623 102 19 96 23 29 31 95 266 105 406 409 OAI222_X1 $T=20950 31800 1 0 $X=20835 $Y=30285
X2624 102 147 96 35 29 31 95 193 379 406 263 OAI222_X1 $T=23800 31800 0 0 $X=23685 $Y=31685
X2625 114 45 96 57 58 59 95 61 385 405 408 OAI222_X1 $T=47740 26200 0 0 $X=47625 $Y=26085
X2626 133 204 96 90 91 65 95 69 365 406 409 OAI222_X1 $T=67880 31800 1 0 $X=67765 $Y=30285
X2628 28 32 95 25 23 96 266 399 406 263 AOI221_X1 $T=19240 31800 1 180 $X=17985 $Y=31685
X2629 330 46 95 290 188 96 64 329 407 408 AOI221_X1 $T=48690 29000 0 180 $X=47435 $Y=27485
X2630 82 51 95 296 67 96 115 297 407 409 AOI221_X1 $T=52490 29000 0 0 $X=52375 $Y=28885
X2631 340 60 95 310 374 96 210 294 405 262 AOI221_X1 $T=63890 26200 0 180 $X=62635 $Y=24685
X2632 365 122 95 311 312 96 128 364 406 409 AOI221_X1 $T=63890 31800 1 0 $X=63775 $Y=30285
X2633 227 185 137 96 397 344 95 406 409 AOI211_X1 $T=6320 31800 1 0 $X=6205 $Y=30285
X2634 185 266 347 96 137 345 95 407 409 AOI211_X1 $T=9740 29000 0 0 $X=9625 $Y=28885
X2635 185 19 348 96 228 269 95 406 409 AOI211_X1 $T=14490 31800 1 0 $X=14375 $Y=30285
X2636 63 64 386 96 334 370 95 406 263 AOI211_X1 $T=49640 31800 0 0 $X=49525 $Y=31685
X2637 67 70 304 96 338 225 95 407 408 AOI211_X1 $T=56290 29000 1 0 $X=56175 $Y=27485
X2638 126 71 389 96 303 388 95 406 263 AOI211_X1 $T=57620 31800 1 180 $X=56555 $Y=31685
X2639 371 56 305 96 306 359 95 406 409 AOI211_X1 $T=58380 31800 1 0 $X=58265 $Y=30285
X2640 400 93 65 96 94 134 95 407 408 AOI211_X1 $T=68450 29000 1 0 $X=68335 $Y=27485
X2641 381 96 95 108 407 408 CLKBUF_X1 $T=27790 29000 0 180 $X=27105 $Y=27485
X2642 43 96 95 40 405 408 CLKBUF_X1 $T=34060 26200 0 0 $X=33945 $Y=26085
X2646 236 237 152 96 197 195 380 381 95 405 408 OAI33_X1 $T=29500 26200 1 180 $X=28055 $Y=26085
X2647 57 285 157 96 112 110 78 384 95 405 408 OAI33_X1 $T=41090 26200 0 0 $X=40975 $Y=26085
X2648 72 91 326 96 163 66 84 387 95 407 408 OAI33_X1 $T=50970 29000 1 0 $X=50855 $Y=27485
X2649 80 298 91 96 133 326 84 296 95 406 409 OAI33_X1 $T=50970 31800 1 0 $X=50855 $Y=30285
X2650 93 298 133 96 91 169 84 334 95 406 263 OAI33_X1 $T=53060 31800 0 0 $X=52945 $Y=31685
X2651 167 326 65 96 90 205 118 362 95 407 409 OAI33_X1 $T=55340 29000 0 0 $X=55225 $Y=28885
X2652 298 167 90 96 204 205 326 168 95 406 263 OAI33_X1 $T=55340 31800 0 0 $X=55225 $Y=31685
X2653 88 167 163 96 118 66 93 301 95 405 408 OAI33_X1 $T=57810 26200 1 180 $X=56365 $Y=26085
X2654 77 218 176 96 170 125 81 310 95 405 262 OAI33_X1 $T=59900 26200 1 0 $X=59785 $Y=24685
X2655 170 167 118 96 308 309 93 306 95 407 409 OAI33_X1 $T=60090 29000 0 0 $X=59975 $Y=28885
X2656 88 84 70 96 92 90 176 175 95 405 262 OAI33_X1 $T=68070 26200 1 0 $X=67955 $Y=24685
X2658 21 141 143 96 95 406 263 NOR2_X2 $T=15820 31800 0 0 $X=15705 $Y=31685
X2659 26 101 319 96 95 407 408 NOR2_X2 $T=20190 29000 0 180 $X=19125 $Y=27485
X2660 378 96 316 271 95 29 407 409 NAND3_X1 $T=20000 29000 1 180 $X=19125 $Y=28885
X2661 375 96 150 151 95 380 405 408 NAND3_X1 $T=27410 26200 0 0 $X=27295 $Y=26085
X2662 287 96 286 48 95 111 406 409 NAND3_X1 $T=42230 31800 0 180 $X=41355 $Y=30285
X2663 286 96 287 115 95 54 407 408 NAND3_X1 $T=42610 29000 1 0 $X=42495 $Y=27485
X2664 325 96 159 49 95 59 405 408 NAND3_X1 $T=43180 26200 0 0 $X=43065 $Y=26085
X2665 117 96 56 57 95 299 407 408 NAND3_X1 $T=46790 29000 1 0 $X=46675 $Y=27485
X2666 165 96 55 161 95 291 406 263 NAND3_X1 $T=46980 31800 0 0 $X=46865 $Y=31685
X2667 184 96 398 165 95 395 405 408 NAND3_X1 $T=49260 26200 0 0 $X=49145 $Y=26085
X2668 232 96 360 297 95 282 405 408 NAND3_X1 $T=51920 26200 1 180 $X=51045 $Y=26085
X2669 84 96 206 207 95 309 405 262 NAND3_X1 $T=57430 26200 1 0 $X=57315 $Y=24685
X2670 73 96 130 61 95 339 405 408 NAND3_X1 $T=58760 26200 0 0 $X=58645 $Y=26085
X2671 392 96 73 174 95 342 405 408 NAND3_X1 $T=68640 26200 1 180 $X=67765 $Y=26085
X2686 396 333 395 329 96 95 295 405 408 AND4_X1 $T=50020 26200 0 0 $X=49905 $Y=26085
X2687 96 18 191 95 99 405 262 XNOR2_X2 $T=15630 26200 0 180 $X=13615 $Y=24685
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 8 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A1 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 9 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_14
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6 7
** N=11 EP=7 IP=0 FDC=10
M0 8 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 11 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 11 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 10 A 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 10 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 9 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 9 B Z 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI21_X2 A VSS B1 ZN B2 VDD 7 8
** N=11 EP=8 IP=0 FDC=12
M0 VSS A 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 A VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN B2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN B1 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 9 B2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 ZN A VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M7 VDD A ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M8 10 B2 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M9 ZN B1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M10 11 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
M11 VDD B2 11 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_15 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 222 223 224 225 226 227 228 229 230 231 232 233 234 235 236 237 238 239 240
+ 241 242 243 244 245 246 247 248 249 250 251 252 253 254 255 256 257 258 259 278
+ 279
** N=467 EP=261 IP=6206 FDC=2074
M0 87 342 76 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=29115 $Y=20690 $D=1
M1 76 342 87 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29305 $Y=20690 $D=1
M2 459 30 76 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29495 $Y=20690 $D=1
M3 342 27 459 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=29685 $Y=20690 $D=1
M4 90 304 76 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=38425 $Y=20690 $D=1
M5 76 304 90 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38615 $Y=20690 $D=1
M6 460 309 76 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38805 $Y=20690 $D=1
M7 90 89 460 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38995 $Y=20690 $D=1
M8 461 89 90 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39185 $Y=20690 $D=1
M9 76 309 461 462 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=39375 $Y=20690 $D=1
M10 87 342 75 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=29115 $Y=21280 $D=0
M11 75 342 87 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29305 $Y=21280 $D=0
M12 342 30 75 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29495 $Y=21280 $D=0
M13 75 27 342 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=29685 $Y=21280 $D=0
M14 75 304 345 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=38425 $Y=21280 $D=0
M15 345 304 75 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38615 $Y=21280 $D=0
M16 90 309 345 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38805 $Y=21280 $D=0
M17 345 89 90 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38995 $Y=21280 $D=0
M18 90 89 345 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39185 $Y=21280 $D=0
M19 345 309 90 465 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=39375 $Y=21280 $D=0
X2275 127 1 76 75 280 464 279 AND2_X1 $T=1000 23400 0 0 $X=885 $Y=23285
X2276 127 2 76 75 334 463 467 AND2_X1 $T=1950 17800 1 0 $X=1835 $Y=16285
X2277 129 284 76 75 281 463 466 AND2_X1 $T=4990 17800 1 180 $X=4115 $Y=17685
X2278 129 283 76 75 445 462 465 AND2_X1 $T=4230 20600 0 0 $X=4115 $Y=20485
X2279 129 285 76 75 282 464 465 AND2_X1 $T=4990 23400 0 180 $X=4115 $Y=21885
X2280 130 6 76 75 372 464 465 AND2_X1 $T=5940 23400 1 0 $X=5825 $Y=21885
X2281 7 177 76 75 286 463 467 AND2_X1 $T=7840 17800 0 180 $X=6965 $Y=16285
X2282 288 286 76 75 375 462 466 AND2_X1 $T=8410 20600 1 0 $X=8295 $Y=19085
X2290 334 3 76 75 5 278 467 DFF_X1 $T=1000 15000 0 0 $X=885 $Y=14885
X2291 281 4 76 75 180 463 466 DFF_X1 $T=4230 17800 1 180 $X=885 $Y=17685
X2292 445 4 76 75 128 462 466 DFF_X1 $T=1000 20600 1 0 $X=885 $Y=19085
X2293 282 4 76 75 126 464 465 DFF_X1 $T=4230 23400 0 180 $X=885 $Y=21885
X2294 280 3 76 75 10 464 279 DFF_X1 $T=1760 23400 0 0 $X=1645 $Y=23285
X2295 372 8 76 75 83 464 465 DFF_X1 $T=6700 23400 1 0 $X=6585 $Y=21885
X2296 218 8 76 75 88 463 467 DFF_X1 $T=29690 17800 1 0 $X=29575 $Y=16285
X2297 219 3 76 75 145 462 466 DFF_X1 $T=32350 20600 1 0 $X=32235 $Y=19085
X2298 33 8 76 75 236 463 466 DFF_X1 $T=35200 17800 0 0 $X=35085 $Y=17685
X2915 454 76 75 425 463 466 INV_X1 $T=6130 17800 0 0 $X=6015 $Y=17685
X2916 427 76 75 283 464 279 INV_X1 $T=7650 23400 1 180 $X=7155 $Y=23285
X2917 177 76 75 414 278 467 INV_X1 $T=7650 15000 0 0 $X=7535 $Y=14885
X2918 182 76 75 285 464 279 INV_X1 $T=7650 23400 0 0 $X=7535 $Y=23285
X2919 428 76 75 284 462 465 INV_X1 $T=9740 20600 1 180 $X=9245 $Y=20485
X2920 79 76 75 287 462 465 INV_X1 $T=11260 20600 1 180 $X=10765 $Y=20485
X2921 296 76 75 378 463 466 INV_X1 $T=13160 17800 1 180 $X=12665 $Y=17685
X2922 14 76 75 80 278 467 INV_X1 $T=13350 15000 0 0 $X=13235 $Y=14885
X2923 81 76 75 384 464 279 INV_X1 $T=15440 23400 0 0 $X=15325 $Y=23285
X2924 132 76 75 430 278 467 INV_X1 $T=15630 15000 0 0 $X=15515 $Y=14885
X2925 13 76 75 446 462 466 INV_X1 $T=16010 20600 1 0 $X=15895 $Y=19085
X2926 134 76 75 385 463 467 INV_X1 $T=16200 17800 1 0 $X=16085 $Y=16285
X2927 16 76 75 386 463 466 INV_X1 $T=17530 17800 1 180 $X=17035 $Y=17685
X2928 387 76 75 431 462 466 INV_X1 $T=18480 20600 1 0 $X=18365 $Y=19085
X2929 188 76 75 294 278 467 INV_X1 $T=19050 15000 0 0 $X=18935 $Y=14885
X2930 447 76 75 391 464 465 INV_X1 $T=20950 23400 0 180 $X=20455 $Y=21885
X2931 295 76 75 394 278 467 INV_X1 $T=20950 15000 0 0 $X=20835 $Y=14885
X2932 18 76 75 15 463 467 INV_X1 $T=22090 17800 0 180 $X=21595 $Y=16285
X2933 436 76 75 297 463 466 INV_X1 $T=22280 17800 1 180 $X=21785 $Y=17685
X2934 191 76 75 226 462 465 INV_X1 $T=23420 20600 0 0 $X=23305 $Y=20485
X2935 341 76 75 173 463 466 INV_X1 $T=26840 17800 0 0 $X=26725 $Y=17685
X2936 12 76 75 194 463 466 INV_X1 $T=27220 17800 0 0 $X=27105 $Y=17685
X2937 434 76 75 32 462 466 INV_X1 $T=27410 20600 1 0 $X=27295 $Y=19085
X2938 172 76 75 84 463 466 INV_X1 $T=27790 17800 0 0 $X=27675 $Y=17685
X2939 300 76 75 421 464 465 INV_X1 $T=28550 23400 1 0 $X=28435 $Y=21885
X2940 197 76 75 38 464 279 INV_X1 $T=37860 23400 0 0 $X=37745 $Y=23285
X2941 34 76 75 35 463 466 INV_X1 $T=40330 17800 1 180 $X=39835 $Y=17685
X2942 438 76 75 36 464 279 INV_X1 $T=40710 23400 1 180 $X=40215 $Y=23285
X2943 51 76 75 42 463 466 INV_X1 $T=41280 17800 0 0 $X=41165 $Y=17685
X2944 45 76 75 50 463 466 INV_X1 $T=42420 17800 0 0 $X=42305 $Y=17685
X2945 311 76 75 94 462 465 INV_X1 $T=42610 20600 0 0 $X=42495 $Y=20485
X2946 52 76 75 57 463 466 INV_X1 $T=45270 17800 1 180 $X=44775 $Y=17685
X2947 349 76 75 350 464 465 INV_X1 $T=44890 23400 1 0 $X=44775 $Y=21885
X2948 44 76 75 97 463 466 INV_X1 $T=45270 17800 0 0 $X=45155 $Y=17685
X2949 315 76 75 149 278 467 INV_X1 $T=46220 15000 1 180 $X=45725 $Y=14885
X2950 39 76 75 357 462 465 INV_X1 $T=48310 20600 0 0 $X=48195 $Y=20485
X2951 49 76 75 43 462 466 INV_X1 $T=49450 20600 0 180 $X=48955 $Y=19085
X2952 113 76 75 125 278 467 INV_X1 $T=52110 15000 0 0 $X=51995 $Y=14885
X2953 153 76 75 159 463 467 INV_X1 $T=52110 17800 1 0 $X=51995 $Y=16285
X2954 319 76 75 405 462 465 INV_X1 $T=52300 20600 0 0 $X=52185 $Y=20485
X2955 106 76 75 60 278 467 INV_X1 $T=55340 15000 1 180 $X=54845 $Y=14885
X2956 326 76 75 363 463 466 INV_X1 $T=55720 17800 1 180 $X=55225 $Y=17685
X2957 212 76 75 406 278 467 INV_X1 $T=57620 15000 1 180 $X=57125 $Y=14885
X2958 107 76 75 73 463 467 INV_X1 $T=57620 17800 1 0 $X=57505 $Y=16285
X2959 61 76 75 111 464 279 INV_X1 $T=58380 23400 1 180 $X=57885 $Y=23285
X2960 407 76 75 162 463 467 INV_X1 $T=58760 17800 0 180 $X=58265 $Y=16285
X2961 328 76 75 115 462 466 INV_X1 $T=61230 20600 1 0 $X=61115 $Y=19085
X2962 410 76 75 66 278 467 INV_X1 $T=62370 15000 0 0 $X=62255 $Y=14885
X2963 370 76 75 329 464 465 INV_X1 $T=63130 23400 1 0 $X=63015 $Y=21885
X2964 47 76 75 118 463 466 INV_X1 $T=64270 17800 0 0 $X=64155 $Y=17685
X2965 117 76 75 330 464 465 INV_X1 $T=64650 23400 0 180 $X=64155 $Y=21885
X2966 56 76 75 53 463 466 INV_X1 $T=65030 17800 1 180 $X=64535 $Y=17685
X2967 119 76 75 424 278 467 INV_X1 $T=65220 15000 1 180 $X=64725 $Y=14885
X2968 74 76 75 72 463 466 INV_X1 $T=65980 17800 1 180 $X=65485 $Y=17685
X2969 411 76 75 120 462 465 INV_X1 $T=66170 20600 0 0 $X=66055 $Y=20485
X2970 109 76 75 167 463 466 INV_X1 $T=66550 17800 0 0 $X=66435 $Y=17685
X2971 105 76 75 70 462 466 INV_X1 $T=67120 20600 1 0 $X=67005 $Y=19085
X2972 54 76 75 122 462 466 INV_X1 $T=68070 20600 0 180 $X=67575 $Y=19085
X2973 371 76 75 332 463 466 INV_X1 $T=68450 17800 1 180 $X=67955 $Y=17685
X2974 116 76 75 69 462 466 INV_X1 $T=68070 20600 1 0 $X=67955 $Y=19085
X3043 241 83 75 9 10 12 76 337 428 464 465 AOI222_X1 $T=9930 23400 1 0 $X=9815 $Y=21885
X3044 241 239 75 9 11 12 76 78 427 464 279 AOI222_X1 $T=9930 23400 0 0 $X=9815 $Y=23285
X3045 241 240 75 9 23 12 76 85 341 464 465 AOI222_X1 $T=22280 23400 1 0 $X=22165 $Y=21885
X3046 87 217 75 300 29 28 76 450 174 464 279 AOI222_X1 $T=29310 23400 1 180 $X=27675 $Y=23285
X3047 417 66 75 424 68 331 76 118 251 463 467 AOI222_X1 $T=63320 17800 1 0 $X=63205 $Y=16285
X3048 119 44 75 71 72 73 76 233 413 278 467 AOI222_X1 $T=66360 15000 0 0 $X=66245 $Y=14885
X3120 12 181 5 76 75 278 467 DLH_X1 $T=6130 15000 1 180 $X=4115 $Y=14885
X3121 12 447 21 76 75 462 466 DLH_X1 $T=23040 20600 0 180 $X=21025 $Y=19085
X3122 12 387 22 76 75 463 467 DLH_X1 $T=22090 17800 1 0 $X=21975 $Y=16285
X3123 12 436 24 76 75 463 466 DLH_X1 $T=22280 17800 0 0 $X=22165 $Y=17685
X3124 12 295 25 76 75 278 467 DLH_X1 $T=23230 15000 0 0 $X=23115 $Y=14885
X3125 28 302 300 76 75 464 465 DLH_X1 $T=31400 23400 1 0 $X=31285 $Y=21885
X3126 28 195 31 76 75 278 467 DLH_X1 $T=33870 15000 1 180 $X=31855 $Y=14885
X3127 90 301 303 76 75 462 465 DLH_X1 $T=31970 20600 0 0 $X=31855 $Y=20485
X3128 28 304 27 76 75 462 465 DLH_X1 $T=35770 20600 1 180 $X=33755 $Y=20485
X3129 90 450 305 76 75 464 465 DLH_X1 $T=35580 23400 1 0 $X=35465 $Y=21885
X3130 90 196 306 76 75 464 279 DLH_X1 $T=35960 23400 0 0 $X=35845 $Y=23285
X3131 90 449 307 76 75 278 467 DLH_X1 $T=36720 15000 0 0 $X=36605 $Y=14885
X3132 134 75 133 387 295 388 76 463 467 NOR4_X1 $T=17340 17800 1 0 $X=17225 $Y=16285
X3133 240 75 253 239 83 433 76 464 279 NOR4_X1 $T=17720 23400 0 0 $X=17605 $Y=23285
X3134 21 75 22 24 25 437 76 463 467 NOR4_X1 $T=25890 17800 1 0 $X=25775 $Y=16285
X3135 344 75 399 96 302 309 76 462 466 NOR4_X1 $T=39000 20600 1 0 $X=38885 $Y=19085
X3136 69 75 105 319 108 404 76 462 465 NOR4_X1 $T=52680 20600 0 0 $X=52565 $Y=20485
X3137 79 76 375 380 184 221 75 462 465 NAND4_X1 $T=12780 20600 0 0 $X=12665 $Y=20485
X3138 388 76 297 136 243 390 75 278 467 NAND4_X1 $T=18100 15000 0 0 $X=17985 $Y=14885
X3139 433 76 138 437 26 395 75 462 465 NAND4_X1 $T=25320 20600 0 0 $X=25205 $Y=20485
X3140 21 76 22 24 25 86 75 463 467 NAND4_X1 $T=27980 17800 1 0 $X=27865 $Y=16285
X3141 203 76 352 204 354 306 75 464 279 NAND4_X1 $T=46030 23400 0 0 $X=45915 $Y=23285
X3142 198 76 38 43 57 150 75 463 466 NAND4_X1 $T=49260 17800 1 180 $X=48195 $Y=17685
X3143 353 76 53 64 102 344 75 463 466 NAND4_X1 $T=52110 17800 1 180 $X=51045 $Y=17685
X3144 157 76 359 104 57 238 75 464 465 NAND4_X1 $T=53440 23400 0 180 $X=52375 $Y=21885
X3145 115 76 330 159 166 210 75 464 465 NAND4_X1 $T=55530 23400 1 0 $X=55415 $Y=21885
X3146 52 75 96 147 76 229 463 467 NOR3_X1 $T=42610 17800 1 0 $X=42495 $Y=16285
X3147 45 75 91 34 76 353 463 466 NOR3_X1 $T=47360 17800 1 180 $X=46485 $Y=17685
X3148 152 75 153 155 76 320 464 465 NOR3_X1 $T=50590 23400 0 180 $X=49715 $Y=21885
X3149 106 75 212 165 76 361 463 467 NOR3_X1 $T=55340 17800 0 180 $X=54465 $Y=16285
X3150 114 75 105 67 76 366 463 466 NOR3_X1 $T=61040 17800 0 0 $X=60925 $Y=17685
X3151 370 75 105 67 76 89 464 279 NOR3_X1 $T=62940 23400 0 0 $X=62825 $Y=23285
X3179 422 47 351 75 350 305 76 464 465 OAI211_X1 $T=46220 23400 0 180 $X=45155 $Y=21885
X3180 443 326 46 75 54 310 76 463 466 OAI211_X1 $T=55720 17800 0 0 $X=55605 $Y=17685
X3181 420 370 409 75 327 321 76 464 279 OAI211_X1 $T=61610 23400 1 180 $X=60545 $Y=23285
X3183 335 287 170 373 76 75 462 465 AOI21_X1 $T=6700 20600 0 0 $X=6585 $Y=20485
X3184 426 7 335 414 76 75 463 466 AOI21_X1 $T=7270 17800 0 0 $X=7155 $Y=17685
X3185 336 288 454 376 76 75 463 467 AOI21_X1 $T=8600 17800 0 180 $X=7725 $Y=16285
X3186 242 14 379 414 76 75 278 467 AOI21_X1 $T=12590 15000 0 0 $X=12475 $Y=14885
X3187 87 421 337 398 76 75 464 465 AOI21_X1 $T=28930 23400 1 0 $X=28815 $Y=21885
X3188 30 301 398 27 76 75 462 465 AOI21_X1 $T=29880 20600 0 0 $X=29765 $Y=20485
X3189 343 36 314 346 76 75 462 465 AOI21_X1 $T=39570 20600 0 0 $X=39455 $Y=20485
X3190 91 38 400 228 76 75 463 467 AOI21_X1 $T=39760 17800 1 0 $X=39645 $Y=16285
X3191 347 311 402 313 76 75 462 466 AOI21_X1 $T=42040 20600 0 180 $X=41165 $Y=19085
X3192 230 44 355 91 76 75 463 467 AOI21_X1 $T=43940 17800 1 0 $X=43825 $Y=16285
X3193 404 60 423 452 76 75 462 465 AOI21_X1 $T=55340 20600 0 0 $X=55225 $Y=20485
X3194 211 65 323 117 76 75 278 467 AOI21_X1 $T=56670 15000 1 180 $X=55795 $Y=14885
X3195 455 423 160 47 76 75 462 465 AOI21_X1 $T=56860 20600 1 180 $X=55985 $Y=20485
X3196 457 62 443 49 76 75 463 466 AOI21_X1 $T=59140 17800 0 0 $X=59025 $Y=17685
X3197 366 63 457 56 76 75 463 467 AOI21_X1 $T=60660 17800 0 180 $X=59785 $Y=16285
X3198 418 70 419 102 76 75 464 465 AOI21_X1 $T=65790 23400 1 0 $X=65675 $Y=21885
X3202 291 288 75 289 290 429 76 463 466 AOI22_X1 $T=9550 17800 0 0 $X=9435 $Y=17685
X3203 379 381 75 80 222 133 76 463 467 AOI22_X1 $T=13160 17800 1 0 $X=13045 $Y=16285
X3204 432 296 75 132 376 385 76 463 466 AOI22_X1 $T=13160 17800 0 0 $X=13045 $Y=17685
X3205 385 132 75 430 296 134 76 463 467 AOI22_X1 $T=15250 17800 1 0 $X=15135 $Y=16285
X3206 84 430 75 385 256 172 76 278 467 AOI22_X1 $T=16010 15000 0 0 $X=15895 $Y=14885
X3207 431 16 75 386 13 387 76 462 466 AOI22_X1 $T=16390 20600 1 0 $X=16275 $Y=19085
X3208 172 431 75 386 137 84 76 463 466 AOI22_X1 $T=19240 17800 1 180 $X=18175 $Y=17685
X3209 172 17 75 135 434 84 76 462 465 AOI22_X1 $T=18860 20600 0 0 $X=18745 $Y=20485
X3210 435 293 75 294 392 295 76 463 466 AOI22_X1 $T=20190 17800 1 180 $X=19125 $Y=17685
X3211 394 188 75 294 293 295 76 463 467 AOI22_X1 $T=20950 17800 0 180 $X=19885 $Y=16285
X3212 297 18 75 15 292 436 76 463 466 AOI22_X1 $T=20950 17800 0 0 $X=20835 $Y=17685
X3213 87 32 75 449 397 28 76 278 467 AOI22_X1 $T=34820 15000 1 180 $X=33755 $Y=14885
X3214 442 230 75 44 401 403 76 462 466 AOI22_X1 $T=43750 20600 1 0 $X=43635 $Y=19085
X3215 232 96 75 44 176 356 76 464 279 AOI22_X1 $T=50020 23400 1 180 $X=48955 $Y=23285
X3216 151 57 75 161 364 111 76 464 279 AOI22_X1 $T=57050 23400 0 0 $X=56935 $Y=23285
X3217 419 155 75 53 420 121 76 464 279 AOI22_X1 $T=65790 23400 0 0 $X=65675 $Y=23285
X3218 235 124 75 234 333 167 76 463 467 AOI22_X1 $T=69400 17800 0 180 $X=68335 $Y=16285
X3219 287 414 76 429 181 136 75 278 467 OAI22_X1 $T=9740 15000 0 0 $X=9625 $Y=14885
X3220 378 392 76 289 132 385 75 463 467 OAI22_X1 $T=12210 17800 1 0 $X=12095 $Y=16285
X3221 389 446 76 338 386 387 75 462 465 OAI22_X1 $T=15440 20600 0 0 $X=15325 $Y=20485
X3222 446 186 76 340 16 431 75 462 465 OAI22_X1 $T=16390 20600 0 0 $X=16275 $Y=20485
X3223 84 394 76 20 294 172 75 278 467 OAI22_X1 $T=21330 15000 0 0 $X=21215 $Y=14885
X3224 84 297 76 189 15 172 75 278 467 OAI22_X1 $T=22280 15000 0 0 $X=22165 $Y=14885
X3225 257 258 76 139 395 140 75 462 466 OAI22_X1 $T=25510 20600 1 0 $X=25395 $Y=19085
X3226 193 21 76 141 194 415 75 278 467 OAI22_X1 $T=26270 15000 0 0 $X=26155 $Y=14885
X3227 355 103 76 148 91 48 75 463 467 OAI22_X1 $T=44700 17800 1 0 $X=44585 $Y=16285
X3228 40 42 76 356 155 47 75 464 465 OAI22_X1 $T=47740 23400 1 0 $X=47625 $Y=21885
X3229 407 233 76 417 214 62 75 278 467 OAI22_X1 $T=63700 15000 1 180 $X=62635 $Y=14885
X3230 54 169 76 371 124 152 75 463 466 OAI22_X1 $T=68450 17800 0 0 $X=68335 $Y=17685
X3231 200 201 76 314 178 75 97 349 464 279 OAI221_X1 $T=43370 23400 0 0 $X=43255 $Y=23285
X3232 355 103 76 46 317 75 319 205 278 467 OAI221_X1 $T=47930 15000 0 0 $X=47815 $Y=14885
X3233 109 234 76 332 74 75 71 331 463 466 OAI221_X1 $T=66930 17800 0 0 $X=66815 $Y=17685
X3234 425 286 374 426 76 75 463 466 OAI21_X1 $T=6510 17800 0 0 $X=6395 $Y=17685
X3235 335 287 373 374 76 75 462 466 OAI21_X1 $T=6510 20600 1 0 $X=6395 $Y=19085
X3236 383 293 223 382 76 75 462 466 OAI21_X1 $T=15250 20600 0 180 $X=14375 $Y=19085
X3237 436 15 383 339 76 75 463 466 OAI21_X1 $T=15250 17800 0 0 $X=15135 $Y=17685
X3238 295 294 432 382 76 75 463 466 OAI21_X1 $T=18290 17800 1 180 $X=17415 $Y=17685
X3239 297 18 435 393 76 75 463 466 OAI21_X1 $T=20190 17800 0 0 $X=20075 $Y=17685
X3240 30 32 415 397 76 75 463 467 OAI21_X1 $T=28930 17800 1 0 $X=28815 $Y=16285
X3241 48 34 416 38 76 75 463 467 OAI21_X1 $T=37860 17800 1 0 $X=37745 $Y=16285
X3242 400 35 346 439 76 75 463 466 OAI21_X1 $T=39950 17800 1 180 $X=39075 $Y=17685
X3243 401 39 303 402 76 75 462 466 OAI21_X1 $T=40520 20600 1 0 $X=40405 $Y=19085
X3244 228 42 347 38 76 75 463 466 OAI21_X1 $T=41660 17800 0 0 $X=41545 $Y=17685
X3245 57 45 403 46 76 75 462 466 OAI21_X1 $T=44700 20600 1 0 $X=44585 $Y=19085
X3246 98 46 316 38 76 75 462 465 OAI21_X1 $T=45650 20600 1 180 $X=44775 $Y=20485
X3247 40 50 318 146 76 75 464 465 OAI21_X1 $T=47740 23400 0 180 $X=46865 $Y=21885
X3248 103 53 324 43 76 75 463 467 OAI21_X1 $T=51350 17800 1 0 $X=51235 $Y=16285
X3249 54 55 101 325 76 75 464 279 OAI21_X1 $T=51730 23400 0 0 $X=51615 $Y=23285
X3250 70 56 441 155 76 75 462 466 OAI21_X1 $T=52110 20600 1 0 $X=51995 $Y=19085
X3251 456 360 442 362 76 75 462 466 OAI21_X1 $T=55150 20600 0 180 $X=54275 $Y=19085
X3252 364 53 408 365 76 75 464 465 OAI21_X1 $T=58570 23400 1 0 $X=58455 $Y=21885
X3253 177 76 77 336 75 278 467 NAND2_X1 $T=8030 15000 0 0 $X=7915 $Y=14885
X3254 376 76 375 426 75 462 466 NAND2_X1 $T=9740 20600 0 180 $X=9055 $Y=19085
X3255 289 76 288 377 75 463 467 NAND2_X1 $T=10310 17800 0 180 $X=9625 $Y=16285
X3256 377 76 7 381 75 463 467 NAND2_X1 $T=10310 17800 1 0 $X=10195 $Y=16285
X3257 136 76 181 288 75 278 467 NAND2_X1 $T=11260 15000 1 180 $X=10575 $Y=14885
X3258 389 76 186 185 75 464 279 NAND2_X1 $T=13350 23400 0 0 $X=13235 $Y=23285
X3259 338 76 292 339 75 462 465 NAND2_X1 $T=14870 20600 1 180 $X=14185 $Y=20485
X3260 383 76 293 382 75 463 466 NAND2_X1 $T=15250 17800 1 180 $X=14565 $Y=17685
X3261 82 76 384 135 75 464 465 NAND2_X1 $T=16960 23400 0 180 $X=16275 $Y=21885
X3262 390 76 391 17 75 464 465 NAND2_X1 $T=19620 23400 0 180 $X=18935 $Y=21885
X3263 340 76 292 393 75 462 465 NAND2_X1 $T=20950 20600 0 0 $X=20835 $Y=20485
X3264 96 76 41 308 75 464 465 NAND2_X1 $T=37480 23400 1 0 $X=37365 $Y=21885
X3265 146 76 38 438 75 464 279 NAND2_X1 $T=38810 23400 1 180 $X=38125 $Y=23285
X3266 146 76 35 311 75 462 466 NAND2_X1 $T=39950 20600 1 0 $X=39835 $Y=19085
X3267 48 76 42 237 75 464 279 NAND2_X1 $T=40710 23400 0 0 $X=40595 $Y=23285
X3268 45 76 42 312 75 464 465 NAND2_X1 $T=42610 23400 0 180 $X=41925 $Y=21885
X3269 94 76 41 348 75 462 465 NAND2_X1 $T=42990 20600 0 0 $X=42875 $Y=20485
X3270 94 76 38 40 75 462 465 NAND2_X1 $T=44320 20600 0 0 $X=44205 $Y=20485
X3271 36 76 34 231 75 463 466 NAND2_X1 $T=47930 17800 1 180 $X=47245 $Y=17685
X3272 357 76 50 153 75 462 465 NAND2_X1 $T=48690 20600 0 0 $X=48575 $Y=20485
X3273 100 76 112 319 75 463 466 NAND2_X1 $T=49830 17800 1 180 $X=49145 $Y=17685
X3274 357 76 46 55 75 462 465 NAND2_X1 $T=49260 20600 0 0 $X=49145 $Y=20485
X3275 100 76 151 152 75 462 466 NAND2_X1 $T=50210 20600 1 0 $X=50095 $Y=19085
X3276 52 76 97 54 75 462 465 NAND2_X1 $T=51160 20600 0 0 $X=51045 $Y=20485
X3277 359 76 405 156 75 464 279 NAND2_X1 $T=53060 23400 1 180 $X=52375 $Y=23285
X3278 363 76 43 322 75 463 467 NAND2_X1 $T=54010 17800 1 0 $X=53895 $Y=16285
X3279 100 76 43 61 75 462 465 NAND2_X1 $T=55340 20600 1 180 $X=54655 $Y=20485
X3280 330 76 65 106 75 464 465 NAND2_X1 $T=55530 23400 0 180 $X=54845 $Y=21885
X3281 104 76 100 328 75 462 466 NAND2_X1 $T=55720 20600 0 180 $X=55035 $Y=19085
X3282 405 76 49 109 75 464 465 NAND2_X1 $T=56480 23400 1 0 $X=56365 $Y=21885
X3283 406 76 165 211 75 278 467 NAND2_X1 $T=57240 15000 1 180 $X=56555 $Y=14885
X3284 104 76 57 110 75 462 465 NAND2_X1 $T=56860 20600 0 0 $X=56745 $Y=20485
X3285 162 76 115 107 75 463 467 NAND2_X1 $T=57620 17800 0 180 $X=56935 $Y=16285
X3286 112 76 97 326 75 463 466 NAND2_X1 $T=58380 17800 1 180 $X=57695 $Y=17685
X3287 359 76 115 164 75 278 467 NAND2_X1 $T=61230 15000 0 0 $X=61115 $Y=14885
X3288 118 76 115 410 75 278 467 NAND2_X1 $T=62370 15000 1 180 $X=61685 $Y=14885
X3289 115 76 56 74 75 463 466 NAND2_X1 $T=61800 17800 0 0 $X=61685 $Y=17685
X3290 116 76 155 369 75 462 466 NAND2_X1 $T=62180 20600 1 0 $X=62065 $Y=19085
X3291 115 76 65 370 75 462 465 NAND2_X1 $T=62370 20600 0 0 $X=62255 $Y=20485
X3292 67 76 53 407 75 463 466 NAND2_X1 $T=63700 17800 0 0 $X=63585 $Y=17685
X3293 330 76 161 62 75 464 279 NAND2_X1 $T=63700 23400 0 0 $X=63585 $Y=23285
X3294 155 76 53 117 75 462 466 NAND2_X1 $T=65410 20600 1 0 $X=65295 $Y=19085
X3295 69 76 70 411 75 462 466 NAND2_X1 $T=65980 20600 1 0 $X=65865 $Y=19085
X3296 122 76 169 444 75 278 467 NAND2_X1 $T=67880 15000 0 0 $X=67765 $Y=14885
X3297 123 76 69 168 75 464 279 NAND2_X1 $T=68640 23400 1 180 $X=67955 $Y=23285
X3298 287 75 414 291 76 462 466 NOR2_X1 $T=10310 20600 0 180 $X=9625 $Y=19085
X3299 82 75 81 187 76 464 279 NOR2_X1 $T=16580 23400 0 0 $X=16465 $Y=23285
X3300 390 75 447 224 76 464 279 NOR2_X1 $T=20380 23400 0 0 $X=20265 $Y=23285
X3301 396 75 448 143 76 462 466 NOR2_X1 $T=27790 20600 1 0 $X=27675 $Y=19085
X3302 348 75 45 92 76 463 467 NOR2_X1 $T=43370 17800 1 0 $X=43255 $Y=16285
X3303 49 75 151 104 76 462 465 NOR2_X1 $T=50590 20600 0 0 $X=50475 $Y=20485
X3304 106 75 207 359 76 464 465 NOR2_X1 $T=54010 23400 0 180 $X=53325 $Y=21885
X3305 59 75 209 158 76 278 467 NOR2_X1 $T=55340 15000 0 0 $X=55225 $Y=14885
X3335 76 378 171 432 75 462 466 XNOR2_X1 $T=11260 20600 1 0 $X=11145 $Y=19085
X3336 76 392 255 296 75 462 466 XNOR2_X1 $T=18860 20600 1 0 $X=18745 $Y=19085
X3337 76 293 248 435 75 462 466 XNOR2_X1 $T=20000 20600 1 0 $X=19885 $Y=19085
X3338 76 192 299 298 75 464 465 XNOR2_X1 $T=24940 23400 1 0 $X=24825 $Y=21885
X3339 76 192 396 27 75 462 465 XNOR2_X1 $T=26270 20600 0 0 $X=26155 $Y=20485
X3340 76 142 27 299 75 464 279 XNOR2_X1 $T=27790 23400 1 180 $X=26535 $Y=23285
X3341 298 19 190 249 75 76 300 464 279 FA_X1 $T=20950 23400 0 0 $X=20835 $Y=23285
X3352 287 77 75 290 291 76 381 131 463 466 AOI221_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X3353 175 144 75 30 31 76 244 227 278 467 AOI221_X1 $T=28740 15000 0 0 $X=28625 $Y=14885
X3354 416 400 75 37 310 76 92 451 278 467 AOI221_X1 $T=39760 15000 0 0 $X=39645 $Y=14885
X3355 308 198 75 40 312 76 41 313 464 465 AOI221_X1 $T=40900 23400 1 0 $X=40785 $Y=21885
X3356 318 51 75 320 321 76 118 354 464 465 AOI221_X1 $T=48690 23400 1 0 $X=48575 $Y=21885
X3357 49 97 75 52 363 76 441 360 463 466 AOI221_X1 $T=52110 17800 0 0 $X=51995 $Y=17685
X3358 323 154 75 324 58 76 60 317 278 467 AOI221_X1 $T=52490 15000 0 0 $X=52375 $Y=14885
X3359 56 57 367 76 151 456 75 462 466 AOI211_X1 $T=57430 20600 0 180 $X=56365 $Y=19085
X3360 369 65 49 76 52 367 75 462 466 AOI211_X1 $T=61230 20600 0 180 $X=60165 $Y=19085
X3361 216 65 328 76 369 368 75 462 465 AOI211_X1 $T=61420 20600 0 0 $X=61305 $Y=20485
X3362 453 329 408 76 368 422 75 464 465 AOI211_X1 $T=63130 23400 0 180 $X=62065 $Y=21885
X3363 412 168 117 76 64 458 75 462 465 AOI211_X1 $T=68450 20600 0 0 $X=68335 $Y=20485
X3368 30 29 76 75 463 466 INV_X2 $T=29690 17800 0 0 $X=29575 $Y=17685
X3369 308 48 34 76 51 50 41 343 75 464 465 OAI33_X1 $T=38050 23400 1 0 $X=37935 $Y=21885
X3370 312 438 112 76 43 201 40 199 75 464 279 OAI33_X1 $T=42040 23400 0 0 $X=41925 $Y=23285
X3371 93 348 50 76 112 202 245 95 75 278 467 OAI33_X1 $T=42800 15000 0 0 $X=42685 $Y=14885
X3372 57 39 45 76 155 47 151 440 75 462 466 OAI33_X1 $T=47740 20600 1 0 $X=47625 $Y=19085
X3373 59 315 52 76 322 358 344 206 75 278 467 OAI33_X1 $T=49070 15000 0 0 $X=48955 $Y=14885
X3374 108 106 325 76 153 107 64 208 75 464 279 OAI33_X1 $T=53060 23400 0 0 $X=52945 $Y=23285
X3375 102 110 407 76 322 62 64 452 75 462 466 OAI33_X1 $T=58950 20600 1 0 $X=58835 $Y=19085
X3376 163 107 153 76 62 410 246 250 75 278 467 OAI33_X1 $T=59900 15000 0 0 $X=59785 $Y=14885
X3377 155 326 49 76 108 411 370 215 75 462 465 OAI33_X1 $T=65410 20600 1 180 $X=63965 $Y=20485
X3378 304 146 302 76 75 462 466 NOR2_X2 $T=35580 20600 1 0 $X=35465 $Y=19085
X3380 17 76 82 384 75 186 464 279 NAND3_X1 $T=16580 23400 1 180 $X=15705 $Y=23285
X3381 135 76 390 391 75 389 464 465 NAND3_X1 $T=18290 23400 1 0 $X=18175 $Y=21885
X3382 416 76 146 51 75 439 463 466 NAND3_X1 $T=38430 17800 0 0 $X=38315 $Y=17685
X3383 406 76 198 38 75 399 462 466 NAND3_X1 $T=42990 20600 1 0 $X=42875 $Y=19085
X3384 48 76 38 259 75 315 278 467 NAND3_X1 $T=46220 15000 0 0 $X=46105 $Y=14885
X3385 316 76 146 91 75 352 464 465 NAND3_X1 $T=46220 23400 1 0 $X=46105 $Y=21885
X3386 440 76 49 97 75 351 462 465 NAND3_X1 $T=47360 20600 1 180 $X=46485 $Y=20485
X3387 99 76 120 65 75 358 463 467 NAND3_X1 $T=49260 17800 1 0 $X=49145 $Y=16285
X3388 361 76 353 363 75 59 463 467 NAND3_X1 $T=54010 17800 0 180 $X=53135 $Y=16285
X3389 405 76 162 105 75 365 462 465 NAND3_X1 $T=58570 20600 0 0 $X=58455 $Y=20485
X3390 209 76 406 102 75 63 278 467 NAND3_X1 $T=59140 15000 0 0 $X=59025 $Y=14885
X3391 111 76 162 116 75 409 464 279 NAND3_X1 $T=59140 23400 0 0 $X=59025 $Y=23285
X3392 114 76 89 157 75 455 462 465 NAND3_X1 $T=59330 20600 0 0 $X=59215 $Y=20485
X3393 213 76 405 330 75 327 464 279 NAND3_X1 $T=59900 23400 0 0 $X=59785 $Y=23285
X3394 247 76 330 329 75 362 464 465 NAND3_X1 $T=64270 23400 0 180 $X=63395 $Y=21885
X3395 330 76 165 70 75 216 464 279 NAND3_X1 $T=65030 23400 0 0 $X=64915 $Y=23285
X3396 406 76 166 53 75 418 462 465 NAND3_X1 $T=66170 20600 1 180 $X=65295 $Y=20485
X3397 102 76 120 166 75 412 462 465 NAND3_X1 $T=67690 20600 0 0 $X=67575 $Y=20485
X3398 444 76 413 333 75 254 278 467 NAND3_X1 $T=68450 15000 0 0 $X=68335 $Y=14885
X3417 293 292 296 13 76 75 380 462 466 AND4_X1 $T=13540 20600 0 180 $X=12285 $Y=19085
X3418 76 13 389 75 183 464 279 XNOR2_X2 $T=11450 23400 0 0 $X=11335 $Y=23285
X3419 207 322 76 75 325 464 465 OR2_X1 $T=52490 23400 0 180 $X=51615 $Y=21885
X3420 458 179 76 75 453 464 465 OR2_X1 $T=68640 23400 1 0 $X=68525 $Y=21885
X3445 75 192 448 142 76 464 465 XOR2_X1 $T=26080 23400 1 0 $X=25965 $Y=21885
X3446 75 252 307 451 76 278 467 XOR2_X1 $T=39760 15000 1 180 $X=38505 $Y=14885
X3447 339 76 292 220 338 75 464 465 OAI21_X2 $T=14110 23400 0 180 $X=12665 $Y=21885
X3448 393 76 292 225 340 75 464 465 OAI21_X2 $T=20950 23400 1 0 $X=20835 $Y=21885
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7 8
** N=14 EP=8 IP=0 FDC=16
M0 13 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 10 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 10 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 14 A 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 11 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 9 A S 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 10 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 12 B VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 10 A 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 11 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT CLKGATETST_X4 SE E CK GCK VSS VDD 7 8
** N=21 EP=8 IP=0 FDC=34
M0 9 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS E 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS 12 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=675 $Y=90 $D=1
M3 18 9 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=865 $Y=90 $D=1
M4 13 12 18 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.555e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=1055 $Y=90 $D=1
M5 19 10 13 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.555e-14 PD=4.6e-07 PS=8.3e-07 $X=1245 $Y=165 $D=1
M6 VSS 11 19 7 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=1435 $Y=165 $D=1
M7 11 13 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=3.58e-14 PD=1.04e-06 PS=1.12e-06 $X=1630 $Y=90 $D=1
M8 VSS CK 12 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=2.31e-14 PD=1.14e-06 PS=6.4e-07 $X=2030 $Y=90 $D=1
M9 20 CK VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=2235 $Y=90 $D=1
M10 14 13 20 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2425 $Y=90 $D=1
M11 21 13 14 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2615 $Y=90 $D=1
M12 VSS CK 21 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M13 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=2995 $Y=90 $D=1
M14 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=3185 $Y=90 $D=1
M15 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=3375 $Y=90 $D=1
M16 VSS 14 GCK 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=3565 $Y=90 $D=1
M17 15 SE 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M18 VDD E 15 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M19 VDD 12 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=675 $Y=920 $D=0
M20 16 9 VDD 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=865 $Y=890 $D=0
M21 13 10 16 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=3.6075e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=1055 $Y=890 $D=0
M22 17 12 13 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.6075e-14 PD=4.6e-07 PS=1.12e-06 $X=1245 $Y=1145 $D=0
M23 VDD 11 17 8 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=1435 $Y=1145 $D=0
M24 11 13 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=5.085e-14 PD=1.47e-06 PS=1.55e-06 $X=1630 $Y=680 $D=0
M25 VDD CK 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=7.5425e-14 AS=4.5675e-14 PD=1.57e-06 PS=9.2e-07 $X=2030 $Y=865 $D=0
M26 14 CK VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=7.5425e-14 PD=1.54e-06 PS=1.57e-06 $X=2235 $Y=680 $D=0
M27 VDD 13 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2425 $Y=680 $D=0
M28 14 13 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2615 $Y=680 $D=0
M29 VDD CK 14 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
M30 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=2995 $Y=680 $D=0
M31 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3185 $Y=680 $D=0
M32 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=3375 $Y=680 $D=0
M33 VDD 14 GCK 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 226 227
** N=390 EP=217 IP=4643 FDC=1896
X1780 68 1 70 69 375 227 389 AND2_X1 $T=1000 6600 0 0 $X=885 $Y=6485
X1781 68 2 70 69 376 387 389 AND2_X1 $T=1000 9400 1 0 $X=885 $Y=7885
X1782 68 3 70 69 338 386 388 AND2_X1 $T=1000 12200 1 0 $X=885 $Y=10685
X1783 68 4 70 69 356 226 390 AND2_X1 $T=2520 15000 0 180 $X=1645 $Y=13485
X1784 145 228 70 69 180 227 389 AND2_X1 $T=6130 6600 0 0 $X=6015 $Y=6485
X1785 145 237 70 69 185 227 389 AND2_X1 $T=24180 6600 0 0 $X=24065 $Y=6485
X1786 145 19 70 69 188 227 389 AND2_X1 $T=29120 6600 0 0 $X=29005 $Y=6485
X1787 169 256 70 69 261 387 388 AND2_X1 $T=54960 9400 0 0 $X=54845 $Y=9285
X1788 287 261 70 69 86 387 388 AND2_X1 $T=56860 9400 0 0 $X=56745 $Y=9285
X1789 120 65 70 69 94 387 388 AND2_X1 $T=64080 9400 0 0 $X=63965 $Y=9285
X1799 338 5 70 69 234 387 388 DFF_X1 $T=1000 9400 0 0 $X=885 $Y=9285
X1800 356 5 70 69 232 386 390 DFF_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X1801 375 5 70 69 229 227 389 DFF_X1 $T=1760 6600 0 0 $X=1645 $Y=6485
X1802 376 5 70 69 230 387 389 DFF_X1 $T=1760 9400 1 0 $X=1645 $Y=7885
X1803 176 11 70 69 150 387 389 DFF_X1 $T=10310 9400 1 0 $X=10195 $Y=7885
X1804 9 5 70 69 235 227 389 DFF_X1 $T=10690 6600 0 0 $X=10575 $Y=6485
X1805 177 11 70 69 13 387 389 DFF_X1 $T=13540 9400 1 0 $X=13425 $Y=7885
X1806 193 5 70 69 236 227 389 DFF_X1 $T=17150 6600 1 180 $X=13805 $Y=6485
X1807 178 11 70 69 160 227 389 DFF_X1 $T=20950 6600 0 0 $X=20835 $Y=6485
X1808 16 11 70 69 161 227 389 DFF_X1 $T=25890 6600 0 0 $X=25775 $Y=6485
X1809 18 11 70 69 194 386 390 DFF_X1 $T=27790 12200 0 0 $X=27675 $Y=12085
X2232 97 70 69 272 387 389 INV_X1 $T=7080 9400 0 180 $X=6585 $Y=7885
X2233 230 70 69 273 387 389 INV_X1 $T=7080 9400 1 0 $X=6965 $Y=7885
X2234 229 70 69 357 227 389 INV_X1 $T=7270 6600 0 0 $X=7155 $Y=6485
X2235 274 70 69 297 226 390 INV_X1 $T=8600 15000 1 0 $X=8485 $Y=13485
X2236 207 70 69 295 226 390 INV_X1 $T=9550 15000 1 0 $X=9435 $Y=13485
X2237 232 70 69 231 387 389 INV_X1 $T=10310 9400 0 180 $X=9815 $Y=7885
X2238 276 70 69 154 386 390 INV_X1 $T=9930 12200 0 0 $X=9815 $Y=12085
X2239 233 70 69 98 386 390 INV_X1 $T=12210 12200 0 0 $X=12095 $Y=12085
X2240 100 70 69 101 226 390 INV_X1 $T=14680 15000 0 180 $X=14185 $Y=13485
X2241 236 70 69 339 387 388 INV_X1 $T=22660 9400 0 0 $X=22545 $Y=9285
X2242 234 70 69 340 387 388 INV_X1 $T=23800 9400 0 0 $X=23685 $Y=9285
X2243 235 70 69 304 387 388 INV_X1 $T=24560 9400 0 0 $X=24445 $Y=9285
X2244 14 70 69 381 387 389 INV_X1 $T=24940 9400 1 0 $X=24825 $Y=7885
X2245 359 70 69 358 386 390 INV_X1 $T=25320 12200 0 0 $X=25205 $Y=12085
X2246 306 70 69 298 386 388 INV_X1 $T=25510 12200 1 0 $X=25395 $Y=10685
X2247 308 70 69 301 387 389 INV_X1 $T=26270 9400 1 0 $X=26155 $Y=7885
X2248 73 70 69 198 226 390 INV_X1 $T=29120 15000 0 180 $X=28625 $Y=13485
X2249 311 70 69 303 387 389 INV_X1 $T=28930 9400 1 0 $X=28815 $Y=7885
X2250 74 70 69 187 226 390 INV_X1 $T=29500 15000 0 180 $X=29005 $Y=13485
X2251 312 70 69 243 387 388 INV_X1 $T=31400 9400 0 0 $X=31285 $Y=9285
X2252 277 70 69 310 386 388 INV_X1 $T=31970 12200 0 180 $X=31475 $Y=10685
X2253 278 70 69 305 387 389 INV_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X2254 279 70 69 314 387 388 INV_X1 $T=35200 9400 1 180 $X=34705 $Y=9285
X2255 280 70 69 363 386 390 INV_X1 $T=44700 12200 1 180 $X=44205 $Y=12085
X2256 281 70 69 78 226 390 INV_X1 $T=46600 15000 0 180 $X=46105 $Y=13485
X2257 253 70 69 254 386 388 INV_X1 $T=46410 12200 1 0 $X=46295 $Y=10685
X2258 137 70 69 81 226 390 INV_X1 $T=47170 15000 1 0 $X=47055 $Y=13485
X2259 108 70 69 48 226 390 INV_X1 $T=48310 15000 1 0 $X=48195 $Y=13485
X2260 319 70 69 41 386 390 INV_X1 $T=49070 12200 1 180 $X=48575 $Y=12085
X2261 370 70 69 84 387 388 INV_X1 $T=50400 9400 0 0 $X=50285 $Y=9285
X2262 83 70 69 349 386 390 INV_X1 $T=50780 12200 1 180 $X=50285 $Y=12085
X2263 351 70 69 352 387 388 INV_X1 $T=54960 9400 1 180 $X=54465 $Y=9285
X2264 171 70 69 263 386 390 INV_X1 $T=58190 12200 0 0 $X=58075 $Y=12085
X2265 385 70 69 289 387 389 INV_X1 $T=58380 9400 1 0 $X=58265 $Y=7885
X2266 332 70 69 140 227 389 INV_X1 $T=62180 6600 0 0 $X=62065 $Y=6485
X2267 46 70 69 141 387 388 INV_X1 $T=62180 9400 0 0 $X=62065 $Y=9285
X2268 354 70 69 262 386 388 INV_X1 $T=62940 12200 0 180 $X=62445 $Y=10685
X2269 174 70 69 265 386 390 INV_X1 $T=62560 12200 0 0 $X=62445 $Y=12085
X2270 64 70 69 293 227 389 INV_X1 $T=64270 6600 0 0 $X=64155 $Y=6485
X2271 95 70 69 268 227 389 INV_X1 $T=66170 6600 1 180 $X=65675 $Y=6485
X2272 125 70 69 192 387 389 INV_X1 $T=65980 9400 1 0 $X=65865 $Y=7885
X2322 26 238 69 239 20 21 70 342 306 386 388 AOI222_X1 $T=30070 12200 1 0 $X=29955 $Y=10685
X2323 26 23 69 240 20 21 70 199 308 227 389 AOI222_X1 $T=32350 6600 1 180 $X=30715 $Y=6485
X2324 26 24 69 25 21 20 70 377 311 227 389 AOI222_X1 $T=34250 6600 0 0 $X=34135 $Y=6485
X2325 26 27 69 244 20 21 70 344 277 386 388 AOI222_X1 $T=36150 12200 0 180 $X=34515 $Y=10685
X2326 26 30 69 245 20 21 70 365 279 387 388 AOI222_X1 $T=38240 9400 1 180 $X=36605 $Y=9285
X2327 26 29 69 246 20 21 70 378 278 227 389 AOI222_X1 $T=39190 6600 0 0 $X=39075 $Y=6485
X2328 134 48 69 49 50 144 70 52 321 227 389 AOI222_X1 $T=53060 6600 0 0 $X=52945 $Y=6485
X2329 213 271 69 270 67 269 70 79 266 386 388 AOI222_X1 $T=67500 12200 0 180 $X=65865 $Y=10685
X2378 99 274 229 70 69 226 390 DLH_X1 $T=5560 15000 1 0 $X=5445 $Y=13485
X2379 99 149 230 70 69 387 388 DLH_X1 $T=8790 9400 1 180 $X=6775 $Y=9285
X2380 99 276 7 70 69 387 388 DLH_X1 $T=8790 9400 0 0 $X=8675 $Y=9285
X2381 99 147 232 70 69 386 388 DLH_X1 $T=9360 12200 1 0 $X=9245 $Y=10685
X2382 99 233 10 70 69 387 388 DLH_X1 $T=10690 9400 0 0 $X=10575 $Y=9285
X2383 99 148 234 70 69 386 390 DLH_X1 $T=12590 12200 0 0 $X=12475 $Y=12085
X2384 99 183 235 70 69 386 388 DLH_X1 $T=16770 12200 0 180 $X=14755 $Y=10685
X2385 99 100 12 70 69 386 388 DLH_X1 $T=16770 12200 1 0 $X=16655 $Y=10685
X2386 99 103 236 70 69 386 390 DLH_X1 $T=18480 12200 0 0 $X=18365 $Y=12085
X2387 99 196 13 70 69 226 390 DLH_X1 $T=18860 15000 1 0 $X=18745 $Y=13485
X2388 99 156 14 70 69 386 390 DLH_X1 $T=20380 12200 0 0 $X=20265 $Y=12085
X2389 21 312 238 70 69 387 388 DLH_X1 $T=31400 9400 1 180 $X=29385 $Y=9285
X2390 106 342 241 70 69 386 388 DLH_X1 $T=32730 12200 1 0 $X=32615 $Y=10685
X2391 106 313 242 70 69 226 390 DLH_X1 $T=32920 15000 1 0 $X=32805 $Y=13485
X2392 21 40 28 70 69 226 390 DLH_X1 $T=39570 15000 0 180 $X=37555 $Y=13485
X2393 21 80 27 70 69 226 390 DLH_X1 $T=39570 15000 1 0 $X=39455 $Y=13485
X2394 21 61 30 70 69 387 388 DLH_X1 $T=40140 9400 0 0 $X=40025 $Y=9285
X2395 21 57 29 70 69 227 389 DLH_X1 $T=40710 6600 0 0 $X=40595 $Y=6485
X2396 106 344 247 70 69 386 390 DLH_X1 $T=40710 12200 0 0 $X=40595 $Y=12085
X2397 106 365 250 70 69 387 388 DLH_X1 $T=44320 9400 0 0 $X=44205 $Y=9285
X2398 106 378 251 70 69 227 389 DLH_X1 $T=44700 6600 0 0 $X=44585 $Y=6485
X2399 232 69 97 229 230 129 70 386 390 NOR4_X1 $T=7080 12200 0 0 $X=6965 $Y=12085
X2400 183 69 103 147 149 296 70 386 390 NOR4_X1 $T=15440 12200 1 180 $X=14375 $Y=12085
X2401 13 69 7 10 12 157 70 386 388 NOR4_X1 $T=21140 12200 1 0 $X=21025 $Y=10685
X2402 234 69 235 14 236 158 70 386 390 NOR4_X1 $T=23230 12200 1 180 $X=22165 $Y=12085
X2403 232 70 97 229 230 215 69 386 388 NAND4_X1 $T=7460 12200 0 180 $X=6395 $Y=10685
X2404 296 70 102 295 297 152 69 226 390 NAND4_X1 $T=15630 15000 1 0 $X=15515 $Y=13485
X2405 234 70 235 14 236 159 69 386 388 NAND4_X1 $T=23040 12200 1 0 $X=22925 $Y=10685
X2406 364 70 363 362 361 247 69 386 390 NAND4_X1 $T=44320 12200 1 180 $X=43255 $Y=12085
X2407 369 70 323 321 371 250 69 227 389 NAND4_X1 $T=50210 6600 0 0 $X=50095 $Y=6485
X2408 120 70 119 374 294 379 69 387 389 NAND4_X1 $T=62180 9400 0 180 $X=61115 $Y=7885
X2409 122 70 334 335 292 191 69 387 389 NAND4_X1 $T=65030 9400 0 180 $X=63965 $Y=7885
X2410 54 69 55 137 70 287 386 390 NOR3_X1 $T=56290 12200 1 180 $X=55415 $Y=12085
X2427 87 108 331 69 262 373 70 387 388 OAI211_X1 $T=58760 9400 0 0 $X=58645 $Y=9285
X2428 66 58 291 69 264 267 70 386 390 OAI211_X1 $T=61040 12200 1 180 $X=59975 $Y=12085
X2429 121 61 57 69 293 333 70 386 388 OAI211_X1 $T=62940 12200 1 0 $X=62825 $Y=10685
X2432 357 6 130 299 70 69 227 389 AOI21_X1 $T=8410 6600 0 0 $X=8295 $Y=6485
X2433 273 6 195 275 70 69 387 389 AOI21_X1 $T=8410 9400 1 0 $X=8295 $Y=7885
X2434 272 6 228 300 70 69 227 389 AOI21_X1 $T=9170 6600 0 0 $X=9055 $Y=6485
X2435 231 6 131 302 70 69 227 389 AOI21_X1 $T=9930 6600 0 0 $X=9815 $Y=6485
X2436 339 6 184 307 70 69 387 389 AOI21_X1 $T=23040 9400 1 0 $X=22925 $Y=7885
X2437 340 6 237 197 70 69 386 388 AOI21_X1 $T=24750 12200 1 0 $X=24635 $Y=10685
X2438 304 6 132 309 70 69 387 388 AOI21_X1 $T=26650 9400 0 0 $X=26535 $Y=9285
X2439 381 6 17 341 70 69 387 389 AOI21_X1 $T=28930 9400 0 180 $X=28055 $Y=7885
X2440 36 33 133 164 70 69 386 390 AOI21_X1 $T=42610 12200 0 0 $X=42495 $Y=12085
X2441 164 35 200 78 70 69 226 390 AOI21_X1 $T=45460 15000 1 0 $X=45345 $Y=13485
X2442 40 80 83 143 70 69 227 389 AOI21_X1 $T=46600 6600 0 0 $X=46485 $Y=6485
X2443 134 44 348 319 70 69 386 388 AOI21_X1 $T=48310 12200 1 0 $X=48195 $Y=10685
X2444 163 42 382 283 70 69 226 390 AOI21_X1 $T=49450 15000 1 0 $X=49335 $Y=13485
X2445 322 46 350 55 70 69 386 390 AOI21_X1 $T=53250 12200 1 180 $X=52375 $Y=12085
X2446 285 85 327 201 70 69 226 390 AOI21_X1 $T=53440 15000 0 180 $X=52565 $Y=13485
X2447 351 51 328 43 70 69 386 388 AOI21_X1 $T=54200 12200 1 0 $X=54085 $Y=10685
X2448 265 52 284 286 70 69 387 389 AOI21_X1 $T=55340 9400 0 180 $X=54465 $Y=7885
X2449 260 51 288 43 70 69 386 388 AOI21_X1 $T=56480 12200 1 0 $X=56365 $Y=10685
X2450 263 89 283 107 70 69 226 390 AOI21_X1 $T=57430 15000 0 180 $X=56555 $Y=13485
X2451 287 51 139 43 70 69 386 390 AOI21_X1 $T=58190 12200 1 180 $X=57315 $Y=12085
X2452 379 57 258 289 70 69 387 389 AOI21_X1 $T=59520 9400 0 180 $X=58645 $Y=7885
X2453 124 263 264 88 70 69 386 390 AOI21_X1 $T=60090 12200 1 180 $X=59215 $Y=12085
X2454 294 59 384 382 70 69 387 389 AOI21_X1 $T=61230 9400 0 180 $X=60355 $Y=7885
X2455 144 60 257 267 70 69 227 389 AOI21_X1 $T=61420 6600 0 0 $X=61305 $Y=6485
X2456 93 63 335 384 70 69 227 389 AOI21_X1 $T=63510 6600 0 0 $X=63395 $Y=6485
X2457 123 66 355 89 70 69 226 390 AOI21_X1 $T=65030 15000 0 180 $X=64155 $Y=13485
X2458 380 266 354 203 70 69 386 390 AOI21_X1 $T=64460 12200 0 0 $X=64345 $Y=12085
X2460 276 295 69 297 181 233 70 226 390 AOI22_X1 $T=9930 15000 1 0 $X=9815 $Y=13485
X2461 101 149 69 151 182 100 70 226 390 AOI22_X1 $T=12780 15000 1 0 $X=12665 $Y=13485
X2462 155 154 69 295 23 153 70 386 390 AOI22_X1 $T=17530 12200 1 180 $X=16465 $Y=12085
X2463 366 367 69 368 369 318 70 387 389 AOI22_X1 $T=48310 9400 1 0 $X=48195 $Y=7885
X2464 282 189 69 80 320 82 70 387 388 AOI22_X1 $T=49450 9400 0 0 $X=49335 $Y=9285
X2465 124 110 69 82 371 140 70 227 389 AOI22_X1 $T=52110 6600 1 180 $X=51045 $Y=6485
X2466 383 84 69 256 323 324 70 387 389 AOI22_X1 $T=51350 9400 1 0 $X=51235 $Y=7885
X2467 83 111 69 255 325 327 70 226 390 AOI22_X1 $T=51730 15000 1 0 $X=51615 $Y=13485
X2468 190 49 69 111 372 110 70 227 389 AOI22_X1 $T=53060 6600 1 180 $X=51995 $Y=6485
X2469 370 352 69 372 324 284 70 387 389 AOI22_X1 $T=52300 9400 1 0 $X=52185 $Y=7885
X2470 333 90 69 173 259 118 70 386 388 AOI22_X1 $T=61800 12200 0 180 $X=60735 $Y=10685
X2471 91 61 69 58 374 50 70 387 388 AOI22_X1 $T=61230 9400 0 0 $X=61115 $Y=9285
X2472 293 48 69 171 294 124 70 387 389 AOI22_X1 $T=65030 9400 1 0 $X=64915 $Y=7885
X2473 204 336 69 337 380 126 70 226 390 AOI22_X1 $T=66550 15000 1 0 $X=66435 $Y=13485
X2474 153 98 70 238 297 155 69 386 390 OAI22_X1 $T=18480 12200 1 180 $X=17415 $Y=12085
X2475 71 12 70 275 15 358 69 387 388 OAI22_X1 $T=19240 9400 0 0 $X=19125 $Y=9285
X2476 71 10 70 299 15 298 69 387 389 OAI22_X1 $T=20380 9400 0 180 $X=19315 $Y=7885
X2477 71 7 70 300 15 301 69 387 389 OAI22_X1 $T=20380 9400 1 0 $X=20265 $Y=7885
X2478 71 13 70 302 15 303 69 387 389 OAI22_X1 $T=22090 9400 1 0 $X=21975 $Y=7885
X2479 71 186 70 307 15 305 69 387 389 OAI22_X1 $T=26270 9400 0 180 $X=25205 $Y=7885
X2480 71 104 70 309 15 310 69 386 388 OAI22_X1 $T=27030 12200 1 0 $X=26915 $Y=10685
X2481 71 161 70 341 15 314 69 387 388 OAI22_X1 $T=27410 9400 0 0 $X=27295 $Y=9285
X2482 107 168 70 317 36 37 69 386 388 OAI22_X1 $T=45460 12200 1 0 $X=45345 $Y=10685
X2483 37 36 70 38 254 69 39 367 387 388 OAI221_X1 $T=46220 9400 0 0 $X=46105 $Y=9285
X2484 288 138 70 258 257 69 57 251 227 389 OAI221_X1 $T=58000 6600 1 180 $X=56745 $Y=6485
X2485 117 46 70 260 259 69 56 330 387 389 OAI221_X1 $T=58380 9400 0 180 $X=57125 $Y=7885
X2486 162 243 241 343 70 69 387 388 OAI21_X1 $T=34820 9400 1 180 $X=33945 $Y=9285
X2487 348 253 282 81 70 69 386 388 OAI21_X1 $T=48310 12200 0 180 $X=47435 $Y=10685
X2488 143 38 368 95 70 69 227 389 OAI21_X1 $T=48880 6600 0 0 $X=48765 $Y=6485
X2489 167 43 361 349 70 69 386 390 OAI21_X1 $T=49640 12200 0 0 $X=49525 $Y=12085
X2490 326 47 318 328 70 69 386 388 OAI21_X1 $T=52490 12200 1 0 $X=52375 $Y=10685
X2491 98 70 274 146 69 226 390 NAND2_X1 $T=7460 15000 1 0 $X=7345 $Y=13485
X2492 233 70 297 8 69 226 390 NAND2_X1 $T=10880 15000 1 0 $X=10765 $Y=13485
X2493 101 70 151 73 69 226 390 NAND2_X1 $T=14300 15000 0 180 $X=13615 $Y=13485
X2494 162 70 243 343 69 387 388 NAND2_X1 $T=33490 9400 0 0 $X=33375 $Y=9285
X2495 36 70 31 163 69 226 390 NAND2_X1 $T=41470 15000 1 0 $X=41355 $Y=13485
X2496 165 70 77 105 69 226 390 NAND2_X1 $T=43560 15000 1 0 $X=43445 $Y=13485
X2497 320 70 61 366 69 227 389 NAND2_X1 $T=47360 6600 0 0 $X=47245 $Y=6485
X2498 35 70 77 319 69 226 390 NAND2_X1 $T=48880 15000 1 0 $X=48765 $Y=13485
X2499 140 70 168 95 69 227 389 NAND2_X1 $T=49640 6600 0 0 $X=49525 $Y=6485
X2500 325 70 109 252 69 386 390 NAND2_X1 $T=51350 12200 1 180 $X=50665 $Y=12085
X2501 349 70 45 322 69 386 390 NAND2_X1 $T=51350 12200 0 0 $X=51235 $Y=12085
X2502 350 70 115 255 69 386 390 NAND2_X1 $T=52490 12200 1 180 $X=51805 $Y=12085
X2503 84 70 114 326 69 387 388 NAND2_X1 $T=52300 9400 0 0 $X=52185 $Y=9285
X2504 329 70 115 285 69 226 390 NAND2_X1 $T=54960 15000 0 180 $X=54275 $Y=13485
X2505 290 70 81 172 69 226 390 NAND2_X1 $T=58950 15000 0 180 $X=58265 $Y=13485
X2506 33 70 38 332 69 227 389 NAND2_X1 $T=59520 6600 0 0 $X=59405 $Y=6485
X2507 117 70 82 331 69 387 389 NAND2_X1 $T=59520 9400 1 0 $X=59405 $Y=7885
X2508 38 70 89 90 69 227 389 NAND2_X1 $T=60090 6600 0 0 $X=59975 $Y=6485
X2509 91 70 38 291 69 386 388 NAND2_X1 $T=60850 12200 0 180 $X=60165 $Y=10685
X2510 105 69 44 256 70 387 388 NOR2_X1 $T=51350 9400 1 180 $X=50665 $Y=9285
X2511 54 69 38 351 70 387 388 NOR2_X1 $T=54010 9400 0 0 $X=53895 $Y=9285
X2533 70 208 242 343 69 386 390 XNOR2_X1 $T=32920 12200 0 0 $X=32805 $Y=12085
X2539 21 313 69 22 26 70 73 359 226 390 AOI221_X1 $T=31590 15000 0 180 $X=30335 $Y=13485
X2540 317 80 69 249 248 70 85 364 387 388 AOI221_X1 $T=44130 9400 1 180 $X=42875 $Y=9285
X2541 352 55 69 53 170 70 210 286 227 389 AOI221_X1 $T=54580 6600 0 0 $X=54465 $Y=6485
X2542 137 57 69 54 55 70 89 260 386 390 AOI221_X1 $T=56290 12200 0 0 $X=56175 $Y=12085
X2543 202 175 69 355 50 70 58 334 226 390 AOI221_X1 $T=64270 15000 0 180 $X=63015 $Y=13485
X2544 64 48 69 267 268 70 63 216 227 389 AOI221_X1 $T=64650 6600 0 0 $X=64535 $Y=6485
X2545 316 32 43 70 80 249 69 386 388 AOI211_X1 $T=42230 12200 1 0 $X=42115 $Y=10685
X2546 252 35 281 70 105 280 69 386 390 AOI211_X1 $T=45650 12200 0 0 $X=45535 $Y=12085
X2547 79 40 41 70 80 253 69 386 390 AOI211_X1 $T=47740 12200 0 0 $X=47625 $Y=12085
X2548 135 44 109 70 105 383 69 386 388 AOI211_X1 $T=50400 12200 1 0 $X=50285 $Y=10685
X2549 138 45 330 70 136 353 69 387 389 AOI211_X1 $T=57240 9400 0 180 $X=56175 $Y=7885
X2550 353 261 373 70 211 385 69 386 388 AOI211_X1 $T=58190 12200 1 0 $X=58075 $Y=10685
X2553 36 91 37 70 69 387 388 NOR2_X2 $T=42040 9400 0 0 $X=41925 $Y=9285
X2555 7 70 10 12 69 72 387 388 NAND3_X1 $T=21330 9400 0 0 $X=21215 $Y=9285
X2556 209 70 36 31 69 316 226 390 NAND3_X1 $T=42800 15000 0 180 $X=41925 $Y=13485
X2557 142 70 164 165 69 362 226 390 NAND3_X1 $T=42800 15000 1 0 $X=42685 $Y=13485
X2558 76 70 32 38 69 370 386 388 NAND3_X1 $T=44700 12200 1 0 $X=44585 $Y=10685
X2559 81 70 36 33 69 281 386 388 NAND3_X1 $T=47550 12200 0 180 $X=46675 $Y=10685
X2560 322 70 112 114 69 113 386 390 NAND3_X1 $T=53250 12200 0 0 $X=53135 $Y=12085
X2561 116 70 121 114 69 329 226 390 NAND3_X1 $T=55720 15000 0 180 $X=54845 $Y=13485
X2562 212 70 62 265 69 292 387 388 NAND3_X1 $T=63320 9400 0 0 $X=63205 $Y=9285
X2563 48 34 70 69 248 386 388 OR2_X1 $T=43180 12200 1 0 $X=43065 $Y=10685
X2564 239 360 238 70 69 74 386 390 HA_X1 $T=31020 12200 0 0 $X=30905 $Y=12085
X2565 240 346 23 70 69 360 227 389 HA_X1 $T=32350 6600 0 0 $X=32235 $Y=6485
X2566 244 28 27 70 69 345 386 390 HA_X1 $T=36340 12200 0 0 $X=36225 $Y=12085
X2567 377 315 24 70 69 346 387 389 HA_X1 $T=36530 9400 1 0 $X=36415 $Y=7885
X2568 245 345 30 70 69 347 387 388 HA_X1 $T=38240 9400 0 0 $X=38125 $Y=9285
X2569 246 347 29 70 69 315 387 389 HA_X1 $T=40330 9400 0 180 $X=38315 $Y=7885
X2570 290 58 57 70 69 92 226 390 HA_X1 $T=61230 15000 1 0 $X=61115 $Y=13485
X2571 336 171 57 70 69 205 386 390 HA_X1 $T=65220 12200 0 0 $X=65105 $Y=12085
X2572 269 95 57 70 69 127 227 389 HA_X1 $T=67500 6600 0 0 $X=67385 $Y=6485
X2573 270 332 57 70 69 128 387 389 HA_X1 $T=67500 9400 1 0 $X=67385 $Y=7885
X2574 271 293 57 70 69 96 386 388 HA_X1 $T=67500 12200 1 0 $X=67385 $Y=10685
X2575 337 61 57 70 69 206 226 390 HA_X1 $T=67500 15000 1 0 $X=67385 $Y=13485
X2576 70 179 214 166 70 69 387 389 CLKGATETST_X4 $T=44510 9400 1 0 $X=44395 $Y=7885
.ENDS
***************************************
.SUBCKT ICV_17
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 125
** N=194 EP=121 IP=2188 FDC=1070
M0 141 34 34 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=48670 $Y=3500 $D=1
M1 34 140 141 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=48860 $Y=3500 $D=1
M2 34 144 142 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=49200 $Y=3500 $D=1
M3 183 141 34 191 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=49390 $Y=3435 $D=1
M4 145 144 183 191 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.0125e-14 AS=3.85e-14 PD=8.7e-07 PS=8.3e-07 $X=49580 $Y=3435 $D=1
M5 184 142 145 191 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.0125e-14 PD=4.6e-07 PS=8.7e-07 $X=49790 $Y=3550 $D=1
M6 34 143 184 191 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=49980 $Y=3550 $D=1
M7 143 145 34 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.58e-14 PD=1.11e-06 PS=1.12e-06 $X=50175 $Y=3295 $D=1
M8 34 145 143 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=50365 $Y=3295 $D=1
M9 34 43 144 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=3.36e-14 PD=1.14e-06 PS=7.4e-07 $X=50760 $Y=3500 $D=1
M10 185 43 34 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=50965 $Y=3295 $D=1
M11 146 145 185 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51155 $Y=3295 $D=1
M12 186 145 146 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51345 $Y=3295 $D=1
M13 34 43 186 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51535 $Y=3295 $D=1
M14 187 43 34 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51725 $Y=3295 $D=1
M15 146 145 187 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51915 $Y=3295 $D=1
M16 188 145 146 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=52105 $Y=3295 $D=1
M17 34 43 188 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=52295 $Y=3295 $D=1
M18 45 146 34 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=52485 $Y=3515 $D=1
M19 34 146 45 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=52675 $Y=3515 $D=1
M20 45 146 34 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=52865 $Y=3515 $D=1
M21 34 146 45 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=53055 $Y=3515 $D=1
M22 45 146 34 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=53245 $Y=3515 $D=1
M23 34 146 45 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=53435 $Y=3515 $D=1
M24 45 146 34 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=53625 $Y=3515 $D=1
M25 34 146 45 191 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=53815 $Y=3515 $D=1
M26 34 150 48 191 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=55905 $Y=3890 $D=1
M27 189 148 34 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=56095 $Y=3890 $D=1
M28 190 149 189 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=56285 $Y=3890 $D=1
M29 150 49 190 191 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=56475 $Y=3890 $D=1
M30 180 34 141 193 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=48670 $Y=2490 $D=0
M31 46 140 180 193 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=48860 $Y=2490 $D=0
M32 46 144 142 193 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=49200 $Y=2490 $D=0
M33 181 141 46 193 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=49390 $Y=2490 $D=0
M34 145 142 181 193 PMOS_VTL L=5e-08 W=4.2e-07 AD=4.245e-14 AS=5.88e-14 PD=1.16e-06 PS=1.12e-06 $X=49580 $Y=2490 $D=0
M35 182 144 145 193 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=4.245e-14 PD=4.6e-07 PS=1.16e-06 $X=49790 $Y=2630 $D=0
M36 46 143 182 193 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=49980 $Y=2630 $D=0
M37 143 145 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=5.085e-14 PD=1.54e-06 PS=1.55e-06 $X=50175 $Y=2490 $D=0
M38 46 145 143 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=50365 $Y=2490 $D=0
M39 46 43 144 193 PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=5.04e-14 PD=1.57e-06 PS=9.5e-07 $X=50760 $Y=2695 $D=0
M40 146 43 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06 PS=1.57e-06 $X=50965 $Y=2490 $D=0
M41 46 145 146 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51155 $Y=2490 $D=0
M42 146 145 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51345 $Y=2490 $D=0
M43 46 43 146 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51535 $Y=2490 $D=0
M44 146 43 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51725 $Y=2490 $D=0
M45 46 145 146 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51915 $Y=2490 $D=0
M46 146 145 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52105 $Y=2490 $D=0
M47 46 43 146 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52295 $Y=2490 $D=0
M48 45 146 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52485 $Y=2490 $D=0
M49 46 146 45 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52675 $Y=2490 $D=0
M50 45 146 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52865 $Y=2490 $D=0
M51 46 146 45 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=53055 $Y=2490 $D=0
M52 45 146 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=53245 $Y=2490 $D=0
M53 46 146 45 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=53435 $Y=2490 $D=0
M54 45 146 46 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=53625 $Y=2490 $D=0
M55 46 146 45 193 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=53815 $Y=2490 $D=0
M56 46 150 48 194 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=55905 $Y=4480 $D=0
M57 150 148 46 194 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=56095 $Y=4795 $D=0
M58 46 149 150 194 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=56285 $Y=4795 $D=0
M59 150 49 46 194 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=56475 $Y=4795 $D=0
X983 36 2 34 46 173 191 194 AND2_X1 $T=6130 3800 1 180 $X=5255 $Y=3685
X984 36 3 34 46 165 191 194 AND2_X1 $T=6130 3800 0 0 $X=6015 $Y=3685
X985 36 4 34 46 174 191 194 AND2_X1 $T=8410 3800 0 0 $X=8295 $Y=3685
X986 38 6 34 46 138 192 193 AND2_X1 $T=10690 1000 1 180 $X=9815 $Y=885
X987 38 7 34 46 175 192 193 AND2_X1 $T=12210 1000 0 0 $X=12095 $Y=885
X988 53 8 34 46 75 191 193 AND2_X1 $T=12210 3800 1 0 $X=12095 $Y=2285
X989 38 9 34 46 178 192 193 AND2_X1 $T=15440 1000 1 180 $X=14565 $Y=885
X990 38 10 34 46 109 191 194 AND2_X1 $T=15250 3800 0 0 $X=15135 $Y=3685
X991 53 11 34 46 92 125 194 AND2_X1 $T=17150 6600 0 180 $X=16275 $Y=5085
X992 38 12 34 46 93 192 193 AND2_X1 $T=17340 1000 0 0 $X=17225 $Y=885
X993 53 14 34 46 166 191 193 AND2_X1 $T=18670 3800 1 0 $X=18555 $Y=2285
X994 38 15 34 46 77 191 193 AND2_X1 $T=21900 3800 0 180 $X=21025 $Y=2285
X995 36 16 34 46 126 191 194 AND2_X1 $T=21710 3800 0 0 $X=21595 $Y=3685
X996 38 17 34 46 167 191 193 AND2_X1 $T=23610 3800 1 0 $X=23495 $Y=2285
X997 38 18 34 46 78 191 193 AND2_X1 $T=25510 3800 1 0 $X=25395 $Y=2285
X998 36 19 34 46 127 191 194 AND2_X1 $T=27220 3800 0 0 $X=27105 $Y=3685
X999 38 20 34 46 79 191 194 AND2_X1 $T=28740 3800 1 180 $X=27865 $Y=3685
X1000 38 21 34 46 128 191 193 AND2_X1 $T=29310 3800 1 0 $X=29195 $Y=2285
X1001 38 22 34 46 41 191 194 AND2_X1 $T=30830 3800 0 0 $X=30715 $Y=3685
X1002 53 23 34 46 94 191 193 AND2_X1 $T=32160 3800 1 0 $X=32045 $Y=2285
X1003 36 24 34 46 176 191 194 AND2_X1 $T=33680 3800 0 0 $X=33565 $Y=3685
X1004 38 25 34 46 96 191 193 AND2_X1 $T=35200 3800 1 0 $X=35085 $Y=2285
X1011 173 1 34 46 35 192 193 DFF_X1 $T=1000 1000 0 0 $X=885 $Y=885
X1012 89 1 34 46 69 191 194 DFF_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X1013 165 1 34 46 70 192 193 DFF_X1 $T=4230 1000 0 0 $X=4115 $Y=885
X1014 138 5 34 46 52 125 194 DFF_X1 $T=7650 6600 1 0 $X=7535 $Y=5085
X1015 174 1 34 46 37 191 193 DFF_X1 $T=7840 3800 1 0 $X=7725 $Y=2285
X1016 175 5 34 46 110 191 194 DFF_X1 $T=9170 3800 0 0 $X=9055 $Y=3685
X1017 178 5 34 46 76 191 193 DFF_X1 $T=16200 3800 0 180 $X=12855 $Y=2285
X1018 166 13 34 46 54 191 194 DFF_X1 $T=16010 3800 0 0 $X=15895 $Y=3685
X1019 126 1 34 46 39 192 193 DFF_X1 $T=20380 1000 0 0 $X=20265 $Y=885
X1020 90 1 34 46 40 192 193 DFF_X1 $T=23610 1000 0 0 $X=23495 $Y=885
X1021 167 5 34 46 111 191 194 DFF_X1 $T=23990 3800 0 0 $X=23875 $Y=3685
X1022 127 1 34 46 80 192 193 DFF_X1 $T=30260 1000 0 0 $X=30145 $Y=885
X1023 128 5 34 46 55 125 194 DFF_X1 $T=31020 6600 1 0 $X=30905 $Y=5085
X1024 91 1 34 46 71 192 193 DFF_X1 $T=33490 1000 0 0 $X=33375 $Y=885
X1025 176 1 34 46 72 192 193 DFF_X1 $T=36720 1000 0 0 $X=36605 $Y=885
X1146 179 34 46 129 191 194 INV_X1 $T=34440 3800 0 0 $X=34325 $Y=3685
X1147 28 34 46 53 191 193 INV_X1 $T=38620 3800 0 180 $X=38125 $Y=2285
X1148 28 34 46 38 192 193 INV_X1 $T=40330 1000 1 180 $X=39835 $Y=885
X1149 28 34 46 36 191 193 INV_X1 $T=41280 3800 0 180 $X=40785 $Y=2285
X1150 29 34 46 58 125 194 INV_X1 $T=46030 6600 0 180 $X=45535 $Y=5085
X1151 30 34 46 59 125 194 INV_X1 $T=46030 6600 1 0 $X=45915 $Y=5085
X1152 60 34 46 113 125 194 INV_X1 $T=46790 6600 0 180 $X=46295 $Y=5085
X1153 139 34 46 131 191 194 INV_X1 $T=47740 3800 0 0 $X=47625 $Y=3685
X1154 153 34 46 65 191 194 INV_X1 $T=50400 3800 1 180 $X=49905 $Y=3685
X1155 62 34 46 44 125 194 INV_X1 $T=51350 6600 1 0 $X=51235 $Y=5085
X1156 47 34 46 147 191 193 INV_X1 $T=54960 3800 1 0 $X=54845 $Y=2285
X1157 115 34 46 148 191 193 INV_X1 $T=55910 3800 1 0 $X=55795 $Y=2285
X1158 84 34 46 49 125 194 INV_X1 $T=56860 6600 0 180 $X=56365 $Y=5085
X1159 66 34 46 64 125 194 INV_X1 $T=60660 6600 0 180 $X=60165 $Y=5085
X1160 152 34 46 103 125 194 INV_X1 $T=62940 6600 1 0 $X=62825 $Y=5085
X1161 158 34 46 134 191 193 INV_X1 $T=63320 3800 1 0 $X=63205 $Y=2285
X1162 160 34 46 136 191 194 INV_X1 $T=65980 3800 1 180 $X=65485 $Y=3685
X1189 97 95 129 34 46 125 194 DLH_X1 $T=36150 6600 0 180 $X=34135 $Y=5085
X1190 98 130 26 34 46 191 194 DLH_X1 $T=38810 3800 1 180 $X=36795 $Y=3685
X1191 98 133 27 34 46 191 194 DLH_X1 $T=38810 3800 0 0 $X=38695 $Y=3685
X1192 97 112 131 34 46 125 194 DLH_X1 $T=40900 6600 1 0 $X=40785 $Y=5085
X1199 168 30 154 46 32 83 34 191 194 OAI211_X1 $T=54770 3800 0 0 $X=54655 $Y=3685
X1208 163 130 179 42 34 46 125 194 AOI21_X1 $T=36150 6600 1 0 $X=36035 $Y=5085
X1209 149 30 62 86 34 46 191 194 AOI21_X1 $T=50970 3800 0 0 $X=50855 $Y=3685
X1210 169 33 163 135 34 46 191 194 AOI21_X1 $T=61040 3800 0 0 $X=60925 $Y=3685
X1211 114 136 135 133 34 46 191 194 AOI21_X1 $T=65600 3800 1 180 $X=64725 $Y=3685
X1212 116 137 160 84 34 46 125 194 AOI21_X1 $T=65980 6600 0 180 $X=65105 $Y=5085
X1214 148 155 46 177 170 147 34 191 193 AOI22_X1 $T=56860 3800 1 0 $X=56745 $Y=2285
X1215 100 84 46 65 101 64 34 125 194 AOI22_X1 $T=56860 6600 1 0 $X=56745 $Y=5085
X1216 104 67 46 103 137 50 34 125 194 AOI22_X1 $T=63320 6600 1 0 $X=63205 $Y=5085
X1217 106 172 46 105 159 171 34 192 193 AOI22_X1 $T=64460 1000 1 180 $X=63395 $Y=885
X1218 137 84 34 51 67 50 46 125 194 OAI22_X1 $T=65220 6600 0 180 $X=64155 $Y=5085
X1219 162 107 34 158 161 68 46 191 193 OAI22_X1 $T=69400 3800 0 180 $X=68335 $Y=2285
X1220 115 157 34 134 47 46 151 169 191 193 OAI221_X1 $T=59330 3800 1 0 $X=59215 $Y=2285
X1221 105 29 168 153 34 46 191 194 OAI21_X1 $T=52490 3800 1 180 $X=51615 $Y=3685
X1222 104 49 102 156 34 46 125 194 OAI21_X1 $T=59710 6600 0 180 $X=58835 $Y=5085
X1223 113 34 58 153 46 191 194 NAND2_X1 $T=50400 3800 0 0 $X=50285 $Y=3685
X1224 168 34 30 154 46 191 194 NAND2_X1 $T=54200 3800 0 0 $X=54085 $Y=3685
X1225 86 34 49 85 46 191 194 NAND2_X1 $T=58190 3800 0 0 $X=58075 $Y=3685
X1226 64 34 58 156 46 191 194 NAND2_X1 $T=58760 3800 0 0 $X=58645 $Y=3685
X1227 64 34 65 87 46 125 194 NAND2_X1 $T=60280 6600 0 180 $X=59595 $Y=5085
X1228 50 34 152 88 46 125 194 NAND2_X1 $T=61230 6600 1 0 $X=61115 $Y=5085
X1229 170 34 159 164 46 192 193 NAND2_X1 $T=62940 1000 0 0 $X=62825 $Y=885
X1230 163 46 130 42 34 191 194 NOR2_X1 $T=36340 3800 0 0 $X=36225 $Y=3685
X1231 149 46 30 86 34 191 194 NOR2_X1 $T=54200 3800 1 180 $X=53515 $Y=3685
X1232 44 148 46 31 73 34 147 81 125 194 AOI221_X1 $T=54010 6600 1 0 $X=53895 $Y=5085
X1233 164 33 46 135 74 34 133 139 191 194 AOI221_X1 $T=61800 3800 0 0 $X=61685 $Y=3685
X1235 57 28 34 46 132 191 193 OR2_X1 $T=42230 3800 0 180 $X=41355 $Y=2285
X1236 57 28 34 46 56 192 193 OR2_X1 $T=42800 1000 1 180 $X=41925 $Y=885
X1237 57 28 34 46 140 192 193 OR2_X1 $T=42800 1000 0 0 $X=42685 $Y=885
X1238 117 60 29 34 46 149 191 194 HA_X1 $T=48120 3800 0 0 $X=48005 $Y=3685
X1239 120 153 30 34 46 61 192 193 HA_X1 $T=53250 1000 1 180 $X=51235 $Y=885
X1240 63 29 30 34 46 82 192 193 HA_X1 $T=53250 1000 0 0 $X=53135 $Y=885
X1241 118 149 30 34 46 152 192 193 HA_X1 $T=55150 1000 0 0 $X=55035 $Y=885
X1242 155 85 133 34 46 157 192 193 HA_X1 $T=57050 1000 0 0 $X=56935 $Y=885
X1243 177 66 133 34 46 151 192 193 HA_X1 $T=61040 1000 0 0 $X=60925 $Y=885
X1244 172 156 133 34 46 161 192 193 HA_X1 $T=65600 1000 0 0 $X=65485 $Y=885
X1245 171 87 133 34 46 162 192 193 HA_X1 $T=67500 1000 0 0 $X=67385 $Y=885
X1246 119 152 84 34 46 108 191 194 HA_X1 $T=67500 3800 0 0 $X=67385 $Y=3685
X1247 34 132 43 99 34 46 125 194 CLKGATETST_X4 $T=47550 6600 1 0 $X=47435 $Y=5085
.ENDS
***************************************
.SUBCKT fpa_with_regisers VSS VDD result[14] result[13] inputA[31] result[12] inputB[13] result[11] inputB[14] inputB[12] inputA[12] inputA[14] inputA[13] inputB[11] inputA[11] inputB[1] inputB[10] inputB[0] inputA[16] inputA[0]
+ inputA[10] inputA[1] inputA[9] inputB[9] inputA[8] inputB[8] inputB[7] inputB[5] inputB[4] inputB[3] inputB[2] inputA[2] inputA[7] result[10] result[9] result[1] inputA[4] inputB[19] OF clk
+ result[29] result[28] result[30] result[27] inputA[28] inputB[24] inputA[29] inputB[26] inputA[30] inputA[27] inputB[25] inputA[20] result[26] inputA[26] inputA[19] inputA[25] result[23] result[24] inputA[23] inputA[24]
+ inputA[18] inputB[18] result[25] result[19] inputA[17] en reset inputB[31] result[31] result[2] result[7] result[4] result[8] result[6] inputA[6] inputB[6] result[0] inputA[3] result[3] result[5]
+ inputA[5] inputA[15] result[17] result[16] result[15] inputB[20] inputB[17] inputB[16] result[18] inputB[15] inputA[21] inputB[21] inputB[28] result[22] result[21] result[20] inputA[22] inputB[22] inputB[30] inputB[29]
+ inputB[23] inputB[27] 695
** N=725 EP=103 IP=1722 FDC=14578
X0 inputB[31] 109 46 290 inputA[31] 95 96 152 21 22 19 inputB[13] inputB[14] 17 inputB[12] 33 inputA[12] inputA[14] 47 57
+ 40 inputA[13] 69 44 45 inputB[11] inputA[11] 50 inputB[1] 302 49 54 706 inputB[10] 68 63 inputB[0] 61 inputA[16] 64
+ inputA[0] inputA[1] inputA[10] inputA[9] inputB[9] 79 inputA[8] 81 inputB[5] inputB[7] inputB[4] inputB[3] inputB[2] inputA[2] inputA[7] inputA[4] VDD VSS 12 593
+ 594 27 104 42 90 97 result[1] 5 7 9 11 13 result[12] 705 23 101 29 34 604 599
+ 70 544 73 80 85 94 102 result[2] 542 25 35 37 43 596 51 59 55 158 76 600
+ result[7] result[4] inputB[8] 590 14 134 696 56 62 result[8] result[9] 92 result[31] result[13] 591 595 18 592 543 30
+ 32 39 214 598 157 77 550 result[14] result[11] result[10] 28 78 4 8 702 597 66 84 601 99
+ 719
+ ICV_6 $T=0 0 0 0 $X=0 $Y=59685
X1 109 114 112 602 115 124 125 123 603 258 122 57 157 108 56 23 592 18 129 25
+ 543 132 30 29 160 34 133 40 599 44 212 606 147 69 45 152 143 150 94 706
+ 151 551 163 162 164 550 80 607 55 68 63 70 79 612 178 180 102 95 46 92
+ inputB[6] 186 64 50 171 96 190 inputA[3] inputA[6] inputA[5] 290 VDD VSS 7 39 27 161 146 149 596
+ 165 153 54 177 78 192 544 182 183 97 99 113 591 5 32 14 128 17 201 22
+ 130 131 140 139 144 43 598 13 168 174 608 166 188 189 101 104 result[3] result[5] 111 4
+ 116 37 127 549 202 204 142 552 155 169 172 611 184 result[0] 62 120 630 136 107 118
+ 119 135 28 33 35 595 173 605 47 145 141 49 51 610 175 600 84 90 590 8
+ 121 126 604 705 21 19 593 594 137 148 216 702 597 167 181 601 result[6] 12 9 696
+ 158 42 66 85 191 76 138 154 609 156 61 170 176 179 185 187 110 11 159 719
+ 720
+ ICV_8 $T=0 0 0 0 $X=0 $Y=51285
X2 114 109 157 200 124 603 257 69 197 14 62 32 132 39 134 604 144 605 621 80
+ 151 212 206 208 606 213 299 162 215 163 149 696 59 158 76 159 550 164 222 178
+ 169 180 226 225 611 176 177 612 238 171 181 186 246 243 625 626 255 249 247 245
+ 251 252 inputA[15] 96 290 VDD VSS 194 107 121 614 5 125 133 617 139 148 152 160 95
+ 168 552 174 223 182 233 242 101 115 112 7 198 17 22 23 130 131 137 551 143
+ 150 207 209 140 210 211 147 161 220 608 165 170 189 104 result[15] 193 195 119 203 40
+ 214 620 230 227 229 239 237 562 123 599 607 610 118 613 110 116 117 602 258 201
+ 549 205 616 141 618 561 219 218 622 166 231 250 253 623 188 248 191 254 result[17] 235
+ 240 37 122 111 127 615 135 138 146 46 142 217 79 228 232 236 241 244 result[16] 126
+ 128 145 185 183 184 192 113 108 172 224 179 234 187 609 175 120 624 199 619 221
+ 721 720
+ ICV_9 $T=0 0 0 0 $X=0 $Y=42840
X3 inputB[20] 109 194 614 262 261 263 198 199 628 265 120 196 14 337 40 632 260 208 200
+ 257 122 618 132 23 147 162 271 163 143 635 37 150 621 620 213 214 215 278 154
+ 286 622 302 299 254 356 308 95 227 287 180 178 222 59 79 282 294 225 312 226
+ 637 inputB[17] 228 297 641 311 239 448 293 242 inputB[16] 229 245 233 101 396 310 247 640 253
+ 318 710 624 317 188 244 237 360 323 320 315 313 232 325 326 568 231 236 250 643
+ 249 290 328 VSS VDD 193 256 7 112 202 133 136 634 211 123 152 108 275 141 279
+ 281 217 218 219 288 182 298 307 300 306 314 319 190 251 90 633 258 195 5 542
+ 17 627 22 201 197 615 206 616 269 551 161 210 209 144 207 272 277 561 280 220
+ 283 305 296 638 303 189 224 309 230 240 329 316 374 711 322 255 241 result[18] 264 268
+ 266 129 273 274 276 284 223 301 709 inputB[15] 295 327 115 613 602 114 267 130 631 203
+ 707 205 212 619 155 259 216 221 292 639 697 246 623 625 324 125 124 630 270 617
+ 235 238 243 626 156 92 642 204 291 285 289 234 562 708 153 321 252 629 636 304
+ 248 721 725
+ ICV_11 $T=0 0 0 0 $X=0 $Y=33040
X4 inputB[19] inputB[21] 225 333 inputA[21] 644 602 283 331 265 267 339 95 287 122 258 343 646 707 342
+ 338 197 208 332 270 645 618 136 162 414 163 633 647 257 143 274 636 284 178 294
+ 354 648 285 709 652 292 282 698 651 654 448 357 242 366 296 360 365 317 327 658
+ 653 378 638 712 329 306 247 312 438 228 233 394 389 398 320 319 322 295 321 311
+ 390 245 229 376 642 393 714 328 239 313 307 244 310 253 VDD VSS 262 266 133 152
+ 40 161 347 271 346 348 634 92 289 363 293 361 364 710 305 650 301 372 374 369
+ 375 460 377 382 380 323 660 231 297 188 241 465 309 3 90 104 261 115 268 630
+ 17 708 204 345 344 269 273 350 277 351 77 349 275 649 358 189 387 367 298 370
+ 303 362 657 373 232 318 316 640 314 396 386 568 326 249 397 391 335 340 352 359
+ 371 661 395 325 337 341 637 237 631 264 336 206 635 278 167 279 280 703 300 304
+ 713 381 659 315 383 385 388 641 324 250 256 129 147 334 442 655 639 384 643 629
+ 276 182 160 368 697 286 628 632 155 281 355 656 392 291 379 353 428 724 725
+ ICV_13 $T=0 0 0 0 $X=0 $Y=24685
X5 inputB[22] inputB[28] 225 290 399 inputA[22] 403 283 95 331 333 287 336 581 417 412 339 413 647 415
+ 669 420 644 422 421 667 355 294 178 347 424 670 431 359 358 303 242 439 371 367
+ 651 435 653 292 712 443 369 652 229 365 649 305 658 307 372 228 387 449 701 385
+ 380 390 678 329 311 582 233 568 310 376 681 463 713 316 VDD VSS 401 334 663 405
+ 406 408 343 155 352 353 182 286 392 189 357 434 436 298 441 360 438 370 674 447
+ 655 396 444 452 253 379 383 315 306 386 388 295 247 462 660 250 676 460 468 389
+ 3 465 244 466 398 result[20] 90 result[21] 101 104 260 664 407 410 342 409 671 288 220 73
+ 699 350 OF 668 709 710 698 673 440 677 448 309 657 450 394 375 231 451 700 381
+ 232 455 456 680 241 236 464 454 583 263 627 163 419 345 423 656 400 368 397 result[22]
+ 402 335 115 337 262 646 340 411 416 346 666 348 160 173 429 354 650 362 364 366
+ 363 672 442 703 675 446 377 378 249 382 453 384 661 512 393 391 648 704 430 114
+ 645 338 199 634 144 349 427 297 715 654 374 373 458 467 325 356 361 659 332 414
+ 92 404 665 425 437 679 395 210 344 457 459 433 341 461 272 432 662 418 445 722
+ 724
+ ICV_15 $T=0 0 0 0 $X=0 $Y=14885
X6 inputB[29] inputB[30] inputB[23] inputB[27] 225 95 471 401 476 473 283 474 666 479 173 684 483 716 419 178
+ 294 427 486 432 488 182 671 670 415 416 358 439 501 441 387 435 367 588 314 433
+ 447 303 297 448 250 454 701 237 688 245 451 718 379 677 253 384 487 505 692 507
+ 492 582 255 509 459 293 465 90 VDD VSS 160 428 424 425 715 438 674 292 445 443
+ 239 444 687 450 502 500 318 691 504 242 458 508 511 494 466 399 665 287 407 404
+ 417 411 420 672 189 398 374 452 496 228 678 449 376 311 310 503 329 506 680 241
+ 589 714 247 694 464 468 583 259 682 472 482 436 497 686 499 360 690 711 495 462
+ 675 493 323 101 400 664 406 581 341 405 408 155 409 163 413 667 351 418 414 422
+ 485 370 440 434 302 446 490 385 498 717 456 396 390 460 477 475 683 489 469 403
+ 663 412 480 481 421 668 484 700 455 693 679 478 669 470 410 699 423 685 437 676
+ 461 369 463 681 467 402 429 673 689 457 512 325 clk 662 510 722 723
+ ICV_16 $T=0 0 0 0 $X=0 $Y=6485
X7 290 682 470 472 283 inputA[28] inputA[29] inputB[24] inputA[30] inputA[20] inputB[26] inputA[27] 225 inputB[25] inputA[19] 480 inputA[26] inputA[25] 482 inputA[23]
+ inputA[24] inputA[18] inputB[18] 483 inputA[17] 486 432 reset 445 492 253 384 502 VSS result[29] 101 result[27] 104 result[26] result[23]
+ 704 485 clk 497 308 VDD 678 499 691 323 589 471 90 479 420 489 en 501 588 433
+ 717 686 688 692 493 504 239 454 result[28] result[30] result[19] result[25] 687 693 476 474 683 684 716 result[24]
+ 498 505 689 487 500 509 508 506 469 481 484 478 475 430 685 431 189 294 299 494
+ 690 503 507 495 250 462 310 512 477 473 421 488 490 511 453 510 450 718 694 496
+ 723
+ ICV_18 $T=0 0 0 0 $X=0 $Y=0
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
