/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Tue Jan  3 13:44:33 2023
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 341491754 */

module datapath(b_mantissa, a_mantissa, o_mantissa);
   input [23:0]b_mantissa;
   input [23:0]a_mantissa;
   output [47:0]o_mantissa;

   HA_X1 i_0 (.A(n_534), .B(n_549), .CO(n_557), .S(n_556));
   FA_X1 i_1 (.A(n_544), .B(n_550), .CI(n_567), .CO(n_573), .S(n_572));
   HA_X1 i_2 (.A(n_560), .B(n_557), .CO(n_575), .S(n_574));
   FA_X1 i_3 (.A(n_585), .B(n_578), .CI(n_592), .CO(n_599), .S(n_598));
   HA_X1 i_4 (.A(n_575), .B(n_573), .CO(n_601), .S(n_600));
   FA_X1 i_5 (.A(n_579), .B(n_593), .CI(n_617), .CO(n_625), .S(n_624));
   FA_X1 i_6 (.A(n_611), .B(n_604), .CI(n_601), .CO(n_627), .S(n_626));
   HA_X1 i_7 (.A(n_624), .B(n_599), .CO(n_629), .S(n_628));
   FA_X1 i_8 (.A(n_612), .B(n_605), .CI(n_618), .CO(n_652), .S(n_651));
   FA_X1 i_9 (.A(n_646), .B(n_639), .CI(n_632), .CO(n_654), .S(n_653));
   FA_X1 i_10 (.A(n_651), .B(n_625), .CI(n_629), .CO(n_656), .S(n_655));
   HA_X1 i_11 (.A(n_627), .B(n_653), .CO(n_658), .S(n_657));
   FA_X1 i_12 (.A(n_633), .B(n_675), .CI(n_668), .CO(n_689), .S(n_688));
   FA_X1 i_13 (.A(n_661), .B(n_652), .CI(n_682), .CO(n_691), .S(n_690));
   FA_X1 i_14 (.A(n_654), .B(n_688), .CI(n_690), .CO(n_693), .S(n_692));
   HA_X1 i_15 (.A(n_658), .B(n_656), .CO(n_695), .S(n_694));
   FA_X1 i_16 (.A(n_669), .B(n_662), .CI(n_683), .CO(n_726), .S(n_725));
   FA_X1 i_17 (.A(n_718), .B(n_712), .CI(n_705), .CO(n_728), .S(n_727));
   FA_X1 i_18 (.A(n_698), .B(n_725), .CI(n_689), .CO(n_730), .S(n_729));
   FA_X1 i_19 (.A(n_691), .B(n_727), .CI(n_729), .CO(n_732), .S(n_731));
   HA_X1 i_20 (.A(n_695), .B(n_693), .CO(n_734), .S(n_733));
   FA_X1 i_21 (.A(n_719), .B(n_758), .CI(n_751), .CO(n_766), .S(n_765));
   FA_X1 i_22 (.A(n_744), .B(n_737), .CI(n_726), .CO(n_768), .S(n_767));
   FA_X1 i_23 (.A(n_304), .B(n_728), .CI(n_730), .CO(n_770), .S(n_769));
   FA_X1 i_24 (.A(n_767), .B(n_765), .CI(n_769), .CO(n_772), .S(n_771));
   HA_X1 i_25 (.A(n_734), .B(n_732), .CO(n_774), .S(n_773));
   FA_X1 i_26 (.A(n_798), .B(n_791), .CI(n_784), .CO(n_814), .S(n_813));
   FA_X1 i_27 (.A(n_777), .B(n_306), .CI(n_805), .CO(n_816), .S(n_815));
   FA_X1 i_28 (.A(n_766), .B(n_768), .CI(n_813), .CO(n_818), .S(n_817));
   FA_X1 i_29 (.A(n_770), .B(n_815), .CI(n_817), .CO(n_820), .S(n_819));
   HA_X1 i_30 (.A(n_772), .B(n_774), .CO(n_822), .S(n_821));
   FA_X1 i_31 (.A(n_806), .B(n_852), .CI(n_555), .CO(n_862), .S(n_861));
   FA_X1 i_32 (.A(n_307), .B(n_616), .CI(n_814), .CO(n_866), .S(n_865));
   FA_X1 i_33 (.A(n_816), .B(n_566), .CI(n_861), .CO(n_868), .S(n_867));
   FA_X1 i_34 (.A(n_865), .B(n_818), .CI(n_820), .CO(n_870), .S(n_869));
   HA_X1 i_35 (.A(n_867), .B(n_822), .CO(n_872), .S(n_871));
   FA_X1 i_36 (.A(n_847), .B(n_840), .CI(n_833), .CO(n_909), .S(n_908));
   FA_X1 i_37 (.A(n_603), .B(n_896), .CI(n_889), .CO(n_913), .S(n_912));
   FA_X1 i_38 (.A(n_882), .B(n_875), .CI(n_908), .CO(n_915), .S(n_914));
   FA_X1 i_39 (.A(n_568), .B(n_862), .CI(n_619), .CO(n_917), .S(n_916));
   FA_X1 i_40 (.A(n_866), .B(n_914), .CI(n_912), .CO(n_919), .S(n_918));
   FA_X1 i_41 (.A(n_916), .B(n_868), .CI(n_918), .CO(n_921), .S(n_920));
   HA_X1 i_42 (.A(n_870), .B(n_872), .CO(n_923), .S(n_922));
   FA_X1 i_43 (.A(n_909), .B(n_954), .CI(n_947), .CO(n_970), .S(n_969));
   FA_X1 i_44 (.A(n_940), .B(n_933), .CI(n_926), .CO(n_972), .S(n_971));
   FA_X1 i_45 (.A(n_913), .B(n_915), .CI(n_971), .CO(n_976), .S(n_975));
   FA_X1 i_46 (.A(n_969), .B(n_917), .CI(n_620), .CO(n_978), .S(n_977));
   FA_X1 i_47 (.A(n_919), .B(n_975), .CI(n_977), .CO(n_980), .S(n_979));
   HA_X1 i_48 (.A(n_921), .B(n_923), .CO(n_982), .S(n_981));
   FA_X1 i_49 (.A(n_948), .B(n_941), .CI(n_934), .CO(n_1027), .S(n_1026));
   FA_X1 i_50 (.A(n_1026), .B(n_972), .CI(n_970), .CO(n_1035), .S(n_1034));
   FA_X1 i_51 (.A(n_880), .B(n_1034), .CI(n_976), .CO(n_1039), .S(n_1038));
   FA_X1 i_52 (.A(n_622), .B(n_978), .CI(n_1038), .CO(n_1041), .S(n_1040));
   HA_X1 i_53 (.A(n_980), .B(n_982), .CO(n_1043), .S(n_1042));
   FA_X1 i_54 (.A(n_993), .B(n_986), .CI(n_1027), .CO(n_1089), .S(n_1088));
   FA_X1 i_55 (.A(n_1020), .B(n_959), .CI(n_1074), .CO(n_1091), .S(n_1090));
   FA_X1 i_56 (.A(n_1067), .B(n_1060), .CI(n_1053), .CO(n_1093), .S(n_1092));
   FA_X1 i_57 (.A(n_1046), .B(n_615), .CI(n_1088), .CO(n_1095), .S(n_1094));
   FA_X1 i_58 (.A(n_1035), .B(n_1092), .CI(n_1090), .CO(n_1099), .S(n_1098));
   FA_X1 i_59 (.A(n_1094), .B(n_881), .CI(n_623), .CO(n_1101), .S(n_1100));
   FA_X1 i_60 (.A(n_1039), .B(n_1098), .CI(n_1100), .CO(n_1103), .S(n_1102));
   HA_X1 i_61 (.A(n_1041), .B(n_1043), .CO(n_1105), .S(n_1104));
   FA_X1 i_62 (.A(n_1047), .B(n_879), .CI(n_1143), .CO(n_1159), .S(n_1158));
   FA_X1 i_63 (.A(n_1136), .B(n_1129), .CI(n_1122), .CO(n_1161), .S(n_1160));
   FA_X1 i_64 (.A(n_1115), .B(n_1108), .CI(n_1089), .CO(n_1163), .S(n_1162));
   FA_X1 i_65 (.A(n_983), .B(n_1150), .CI(n_1093), .CO(n_1165), .S(n_1164));
   FA_X1 i_66 (.A(n_1091), .B(n_1158), .CI(n_884), .CO(n_1167), .S(n_1166));
   FA_X1 i_67 (.A(n_1095), .B(n_1162), .CI(n_1160), .CO(n_1169), .S(n_1168));
   FA_X1 i_68 (.A(n_1164), .B(n_1099), .CI(n_1166), .CO(n_1171), .S(n_1170));
   FA_X1 i_69 (.A(n_1101), .B(n_1168), .CI(n_1170), .CO(n_1173), .S(n_1172));
   HA_X1 i_70 (.A(n_1103), .B(n_1172), .CO(n_1175), .S(n_1174));
   FA_X1 i_71 (.A(n_1137), .B(n_1130), .CI(n_1123), .CO(n_1227), .S(n_1226));
   FA_X1 i_72 (.A(n_1151), .B(n_1219), .CI(n_1029), .CO(n_1231), .S(n_1230));
   FA_X1 i_73 (.A(n_1226), .B(n_1161), .CI(n_1159), .CO(n_1237), .S(n_1236));
   FA_X1 i_74 (.A(n_1163), .B(n_1165), .CI(n_987), .CO(n_1239), .S(n_1238));
   FA_X1 i_75 (.A(n_1064), .B(n_1230), .CI(n_1167), .CO(n_1241), .S(n_1240));
   FA_X1 i_76 (.A(n_1236), .B(n_1169), .CI(n_1238), .CO(n_1243), .S(n_1242));
   FA_X1 i_77 (.A(n_1240), .B(n_1171), .CI(n_1242), .CO(n_1245), .S(n_1244));
   HA_X1 i_78 (.A(n_1173), .B(n_1244), .CO(n_1247), .S(n_1246));
   FA_X1 i_79 (.A(n_1214), .B(n_1207), .CI(n_1200), .CO(n_1298), .S(n_1297));
   FA_X1 i_80 (.A(n_1227), .B(n_1220), .CI(n_1138), .CO(n_1302), .S(n_1301));
   FA_X1 i_81 (.A(n_1285), .B(n_1278), .CI(n_1271), .CO(n_1304), .S(n_1303));
   FA_X1 i_82 (.A(n_1264), .B(n_1257), .CI(n_1250), .CO(n_1306), .S(n_1305));
   FA_X1 i_83 (.A(n_984), .B(n_1203), .CI(n_1297), .CO(n_1308), .S(n_1307));
   FA_X1 i_84 (.A(n_1069), .B(n_1231), .CI(n_1301), .CO(n_1310), .S(n_1309));
   FA_X1 i_85 (.A(n_1237), .B(n_988), .CI(n_1305), .CO(n_1312), .S(n_1311));
   FA_X1 i_86 (.A(n_1303), .B(n_1309), .CI(n_1307), .CO(n_1314), .S(n_1313));
   FA_X1 i_87 (.A(n_1239), .B(n_1241), .CI(n_1311), .CO(n_1316), .S(n_1315));
   FA_X1 i_88 (.A(n_1243), .B(n_1313), .CI(n_1315), .CO(n_1318), .S(n_1317));
   HA_X1 i_89 (.A(n_1245), .B(n_1247), .CO(n_1320), .S(n_1319));
   FA_X1 i_90 (.A(n_1279), .B(n_1272), .CI(n_1265), .CO(n_1379), .S(n_1378));
   FA_X1 i_91 (.A(n_1298), .B(n_1365), .CI(n_1358), .CO(n_1383), .S(n_1382));
   FA_X1 i_92 (.A(n_1351), .B(n_1344), .CI(n_1337), .CO(n_1385), .S(n_1384));
   FA_X1 i_93 (.A(n_1330), .B(n_1323), .CI(n_1204), .CO(n_1387), .S(n_1386));
   FA_X1 i_94 (.A(n_1378), .B(n_1372), .CI(n_1306), .CO(n_1389), .S(n_1388));
   FA_X1 i_95 (.A(n_1304), .B(n_1302), .CI(n_1308), .CO(n_1391), .S(n_1390));
   FA_X1 i_96 (.A(n_1386), .B(n_1384), .CI(n_1382), .CO(n_1393), .S(n_1392));
   FA_X1 i_97 (.A(n_1310), .B(n_1390), .CI(n_1388), .CO(n_1395), .S(n_1394));
   FA_X1 i_98 (.A(n_1312), .B(n_1314), .CI(n_1392), .CO(n_1397), .S(n_1396));
   FA_X1 i_99 (.A(n_1316), .B(n_1394), .CI(n_1396), .CO(n_1399), .S(n_1398));
   HA_X1 i_100 (.A(n_1318), .B(n_1398), .CO(n_1401), .S(n_1400));
   FA_X1 i_101 (.A(n_1359), .B(n_1352), .CI(n_1345), .CO(n_1460), .S(n_1459));
   FA_X1 i_102 (.A(n_1379), .B(n_1373), .CI(n_1452), .CO(n_1464), .S(n_1463));
   FA_X1 i_103 (.A(n_1459), .B(n_1385), .CI(n_1383), .CO(n_1472), .S(n_1471));
   FA_X1 i_104 (.A(n_1463), .B(n_1389), .CI(n_1387), .CO(n_1474), .S(n_1473));
   FA_X1 i_105 (.A(n_1391), .B(n_1471), .CI(n_1393), .CO(n_1478), .S(n_1477));
   FA_X1 i_106 (.A(n_1473), .B(n_1395), .CI(n_1209), .CO(n_1480), .S(n_1479));
   FA_X1 i_107 (.A(n_1477), .B(n_1397), .CI(n_1479), .CO(n_1482), .S(n_1481));
   HA_X1 i_108 (.A(n_1399), .B(n_1481), .CO(n_1484), .S(n_1483));
   FA_X1 i_109 (.A(n_1447), .B(n_1440), .CI(n_1433), .CO(n_1544), .S(n_1543));
   FA_X1 i_110 (.A(n_1426), .B(n_1419), .CI(n_1412), .CO(n_1546), .S(n_1545));
   FA_X1 i_111 (.A(n_1405), .B(n_1205), .CI(n_1460), .CO(n_1548), .S(n_1547));
   FA_X1 i_112 (.A(n_1453), .B(n_1536), .CI(n_1530), .CO(n_1550), .S(n_1549));
   FA_X1 i_113 (.A(n_1523), .B(n_1516), .CI(n_1509), .CO(n_1552), .S(n_1551));
   FA_X1 i_114 (.A(n_1502), .B(n_1495), .CI(n_1486), .CO(n_1554), .S(n_1553));
   FA_X1 i_115 (.A(n_1545), .B(n_1543), .CI(n_1201), .CO(n_1556), .S(n_1555));
   FA_X1 i_116 (.A(n_1202), .B(n_1464), .CI(n_1547), .CO(n_1558), .S(n_1557));
   FA_X1 i_117 (.A(n_1472), .B(n_1208), .CI(n_1553), .CO(n_1560), .S(n_1559));
   FA_X1 i_118 (.A(n_1551), .B(n_1549), .CI(n_1474), .CO(n_1562), .S(n_1561));
   FA_X1 i_119 (.A(n_1557), .B(n_1555), .CI(n_1210), .CO(n_1564), .S(n_1563));
   FA_X1 i_120 (.A(n_1559), .B(n_1478), .CI(n_1561), .CO(n_1566), .S(n_1565));
   FA_X1 i_121 (.A(n_1563), .B(n_1480), .CI(n_1565), .CO(n_1568), .S(n_1567));
   HA_X1 i_122 (.A(n_1482), .B(n_1567), .CO(n_1570), .S(n_1569));
   FA_X1 i_123 (.A(n_1510), .B(n_1503), .CI(n_1496), .CO(n_1632), .S(n_1631));
   FA_X1 i_124 (.A(n_1487), .B(n_1546), .CI(n_1544), .CO(n_1634), .S(n_1633));
   FA_X1 i_125 (.A(n_1416), .B(n_1572), .CI(n_1548), .CO(n_1640), .S(n_1639));
   FA_X1 i_126 (.A(n_1631), .B(n_1434), .CI(n_1554), .CO(n_1642), .S(n_1641));
   FA_X1 i_127 (.A(n_1552), .B(n_1550), .CI(n_1633), .CO(n_1644), .S(n_1643));
   FA_X1 i_128 (.A(n_1556), .B(n_1639), .CI(n_1438), .CO(n_1646), .S(n_1645));
   FA_X1 i_129 (.A(n_1441), .B(n_1558), .CI(n_1643), .CO(n_1648), .S(n_1647));
   FA_X1 i_130 (.A(n_1641), .B(n_1560), .CI(n_1562), .CO(n_1650), .S(n_1649));
   FA_X1 i_131 (.A(n_1564), .B(n_1645), .CI(n_1647), .CO(n_1652), .S(n_1651));
   FA_X1 i_132 (.A(n_1649), .B(n_1566), .CI(n_1651), .CO(n_1654), .S(n_1653));
   HA_X1 i_133 (.A(n_1568), .B(n_1653), .CO(n_1656), .S(n_1655));
   FA_X1 i_134 (.A(n_1582), .B(n_1573), .CI(n_1632), .CO(n_1712), .S(n_1711));
   FA_X1 i_135 (.A(n_1695), .B(n_1688), .CI(n_1681), .CO(n_1716), .S(n_1715));
   FA_X1 i_136 (.A(n_1674), .B(n_1667), .CI(n_1658), .CO(n_1718), .S(n_1717));
   FA_X1 i_137 (.A(n_1634), .B(n_1711), .CI(n_1436), .CO(n_1720), .S(n_1719));
   FA_X1 i_138 (.A(n_1640), .B(n_1435), .CI(n_1642), .CO(n_1724), .S(n_1723));
   FA_X1 i_139 (.A(n_1717), .B(n_1715), .CI(n_1644), .CO(n_1726), .S(n_1725));
   FA_X1 i_140 (.A(n_1442), .B(n_1719), .CI(n_1646), .CO(n_1728), .S(n_1727));
   FA_X1 i_141 (.A(n_1723), .B(n_1648), .CI(n_1650), .CO(n_1730), .S(n_1729));
   FA_X1 i_142 (.A(n_1725), .B(n_1727), .CI(n_1652), .CO(n_1732), .S(n_1731));
   FA_X1 i_143 (.A(n_1729), .B(n_1731), .CI(n_1654), .CO(n_1734), .S(n_1733));
   FA_X1 i_144 (.A(n_1703), .B(n_1696), .CI(n_1689), .CO(n_1787), .S(n_1786));
   FA_X1 i_145 (.A(n_1682), .B(n_1675), .CI(n_1668), .CO(n_1789), .S(n_1788));
   FA_X1 i_146 (.A(n_1779), .B(n_1773), .CI(n_1766), .CO(n_1793), .S(n_1792));
   FA_X1 i_147 (.A(n_1759), .B(n_1752), .CI(n_1745), .CO(n_1795), .S(n_1794));
   FA_X1 i_148 (.A(n_1736), .B(n_1712), .CI(n_1788), .CO(n_1797), .S(n_1796));
   FA_X1 i_149 (.A(n_1786), .B(n_1718), .CI(n_1716), .CO(n_1799), .S(n_1798));
   FA_X1 i_150 (.A(n_1720), .B(n_1794), .CI(n_1792), .CO(n_1803), .S(n_1802));
   FA_X1 i_151 (.A(n_1796), .B(n_1724), .CI(n_1798), .CO(n_1805), .S(n_1804));
   FA_X1 i_152 (.A(n_1726), .B(n_1443), .CI(n_1728), .CO(n_1807), .S(n_1806));
   FA_X1 i_153 (.A(n_1802), .B(n_1804), .CI(n_1730), .CO(n_1809), .S(n_1808));
   FA_X1 i_154 (.A(n_1806), .B(n_1732), .CI(n_1808), .CO(n_1811), .S(n_1810));
   FA_X1 i_155 (.A(n_1774), .B(n_1767), .CI(n_1760), .CO(n_1864), .S(n_1863));
   FA_X1 i_156 (.A(n_1753), .B(n_1746), .CI(n_1737), .CO(n_1866), .S(n_1865));
   FA_X1 i_157 (.A(n_1789), .B(n_1787), .CI(n_1857), .CO(n_1868), .S(n_1867));
   FA_X1 i_158 (.A(n_1850), .B(n_1843), .CI(n_1836), .CO(n_1870), .S(n_1869));
   FA_X1 i_159 (.A(n_1437), .B(n_1865), .CI(n_1863), .CO(n_1874), .S(n_1873));
   FA_X1 i_160 (.A(n_1795), .B(n_1793), .CI(n_1867), .CO(n_1876), .S(n_1875));
   FA_X1 i_161 (.A(n_1799), .B(n_1797), .CI(n_1612), .CO(n_1878), .S(n_1877));
   FA_X1 i_162 (.A(n_1869), .B(n_1444), .CI(n_1875), .CO(n_1880), .S(n_1879));
   FA_X1 i_163 (.A(n_1873), .B(n_1803), .CI(n_1877), .CO(n_1882), .S(n_1881));
   FA_X1 i_164 (.A(n_1805), .B(n_1879), .CI(n_1807), .CO(n_1884), .S(n_1883));
   FA_X1 i_165 (.A(n_1881), .B(n_1809), .CI(n_1883), .CO(n_1886), .S(n_1885));
   FA_X1 i_166 (.A(b_mantissa[5]), .B(n_1851), .CI(n_1844), .CO(n_1931), 
      .S(n_1930));
   FA_X1 i_167 (.A(n_1837), .B(n_1830), .CI(n_1823), .CO(n_1933), .S(n_1932));
   FA_X1 i_168 (.A(n_1814), .B(n_1866), .CI(n_1864), .CO(n_1935), .S(n_1934));
   FA_X1 i_169 (.A(n_1858), .B(n_1925), .CI(n_1918), .CO(n_1937), .S(n_1936));
   FA_X1 i_170 (.A(n_1888), .B(n_1932), .CI(n_1930), .CO(n_1941), .S(n_1940));
   FA_X1 i_171 (.A(n_1613), .B(n_1870), .CI(n_1868), .CO(n_1943), .S(n_1942));
   FA_X1 i_172 (.A(n_1934), .B(n_1874), .CI(n_1666), .CO(n_1945), .S(n_1944));
   FA_X1 i_173 (.A(n_1936), .B(n_1876), .CI(n_1942), .CO(n_1947), .S(n_1946));
   FA_X1 i_174 (.A(n_1940), .B(n_1878), .CI(n_1944), .CO(n_1949), .S(n_1948));
   FA_X1 i_175 (.A(n_1880), .B(n_1946), .CI(n_1882), .CO(n_1951), .S(n_1950));
   FA_X1 i_176 (.A(n_1948), .B(n_1884), .CI(n_1950), .CO(n_1953), .S(n_1952));
   FA_X1 i_177 (.A(n_1933), .B(n_1931), .CI(n_1991), .CO(n_2003), .S(n_2002));
   FA_X1 i_178 (.A(n_1985), .B(n_1978), .CI(n_1971), .CO(n_2005), .S(n_2004));
   FA_X1 i_179 (.A(n_1964), .B(n_1955), .CI(n_1935), .CO(n_2007), .S(n_2006));
   FA_X1 i_180 (.A(n_1937), .B(n_2002), .CI(n_1943), .CO(n_2011), .S(n_2010));
   FA_X1 i_181 (.A(n_1941), .B(n_2006), .CI(n_2004), .CO(n_2013), .S(n_2012));
   FA_X1 i_182 (.A(n_1669), .B(n_1945), .CI(n_2010), .CO(n_2015), .S(n_2014));
   FA_X1 i_183 (.A(n_1947), .B(n_2012), .CI(n_1949), .CO(n_2017), .S(n_2016));
   FA_X1 i_184 (.A(n_2014), .B(n_1951), .CI(n_2016), .CO(n_2019), .S(n_2018));
   FA_X1 i_185 (.A(n_1986), .B(n_1979), .CI(n_1972), .CO(n_2065), .S(n_2064));
   FA_X1 i_186 (.A(n_1965), .B(n_1956), .CI(n_1664), .CO(n_2067), .S(n_2066));
   FA_X1 i_187 (.A(n_1665), .B(n_2058), .CI(n_2051), .CO(n_2069), .S(n_2068));
   FA_X1 i_188 (.A(n_2044), .B(n_2037), .CI(n_2030), .CO(n_2071), .S(n_2070));
   FA_X1 i_189 (.A(n_2021), .B(n_2066), .CI(n_2064), .CO(n_2073), .S(n_2072));
   FA_X1 i_190 (.A(n_2005), .B(n_2003), .CI(n_2007), .CO(n_2075), .S(n_2074));
   FA_X1 i_191 (.A(n_1670), .B(n_2070), .CI(n_2068), .CO(n_2077), .S(n_2076));
   FA_X1 i_192 (.A(n_2011), .B(n_2074), .CI(n_2072), .CO(n_2079), .S(n_2078));
   FA_X1 i_193 (.A(n_2013), .B(n_2076), .CI(n_2015), .CO(n_2081), .S(n_2080));
   FA_X1 i_194 (.A(n_2078), .B(n_2017), .CI(n_2080), .CO(n_2083), .S(n_2082));
   FA_X1 i_195 (.A(b_mantissa[8]), .B(n_2052), .CI(n_2045), .CO(n_1), .S(n_0));
   FA_X1 i_196 (.A(n_2038), .B(n_2031), .CI(n_2022), .CO(n_3), .S(n_2));
   FA_X1 i_197 (.A(n_2065), .B(n_2059), .CI(n_265), .CO(n_5), .S(n_4));
   FA_X1 i_198 (.A(n_2108), .B(n_2101), .CI(n_2094), .CO(n_7), .S(n_6));
   FA_X1 i_199 (.A(n_2085), .B(n_2067), .CI(n_2), .CO(n_9), .S(n_8));
   FA_X1 i_200 (.A(n_0), .B(n_2071), .CI(n_2069), .CO(n_11), .S(n_10));
   FA_X1 i_201 (.A(n_4), .B(n_2073), .CI(n_2075), .CO(n_13), .S(n_12));
   FA_X1 i_202 (.A(n_6), .B(n_8), .CI(n_10), .CO(n_15), .S(n_14));
   FA_X1 i_203 (.A(n_2077), .B(n_12), .CI(n_2079), .CO(n_17), .S(n_16));
   FA_X1 i_204 (.A(n_14), .B(n_2081), .CI(n_16), .CO(n_19), .S(n_18));
   FA_X1 i_205 (.A(n_264), .B(n_2109), .CI(n_2102), .CO(n_21), .S(n_20));
   FA_X1 i_206 (.A(n_2095), .B(n_2086), .CI(n_3), .CO(n_23), .S(n_22));
   FA_X1 i_207 (.A(n_1), .B(n_263), .CI(n_262), .CO(n_25), .S(n_24));
   FA_X1 i_208 (.A(n_261), .B(n_260), .CI(n_259), .CO(n_27), .S(n_26));
   FA_X1 i_209 (.A(n_22), .B(n_20), .CI(n_7), .CO(n_29), .S(n_28));
   FA_X1 i_210 (.A(n_5), .B(n_11), .CI(n_9), .CO(n_31), .S(n_30));
   FA_X1 i_211 (.A(n_26), .B(n_24), .CI(n_13), .CO(n_33), .S(n_32));
   FA_X1 i_212 (.A(n_28), .B(n_30), .CI(n_15), .CO(n_35), .S(n_34));
   FA_X1 i_213 (.A(n_32), .B(n_17), .CI(n_34), .CO(n_37), .S(n_36));
   FA_X1 i_214 (.A(n_258), .B(n_256), .CI(n_255), .CO(n_39), .S(n_38));
   FA_X1 i_215 (.A(n_247), .B(n_21), .CI(n_246), .CO(n_41), .S(n_40));
   FA_X1 i_216 (.A(n_245), .B(n_244), .CI(n_243), .CO(n_43), .S(n_42));
   FA_X1 i_217 (.A(n_242), .B(n_23), .CI(n_38), .CO(n_45), .S(n_44));
   FA_X1 i_218 (.A(n_27), .B(n_25), .CI(n_40), .CO(n_47), .S(n_46));
   FA_X1 i_219 (.A(n_29), .B(n_42), .CI(n_44), .CO(n_49), .S(n_48));
   FA_X1 i_220 (.A(n_31), .B(n_46), .CI(n_33), .CO(n_51), .S(n_50));
   FA_X1 i_221 (.A(n_48), .B(n_35), .CI(n_50), .CO(n_53), .S(n_52));
   FA_X1 i_222 (.A(b_mantissa[11]), .B(n_241), .CI(n_240), .CO(n_55), .S(n_54));
   FA_X1 i_223 (.A(n_239), .B(n_238), .CI(n_39), .CO(n_57), .S(n_56));
   FA_X1 i_224 (.A(n_237), .B(n_236), .CI(n_235), .CO(n_59), .S(n_58));
   FA_X1 i_225 (.A(n_234), .B(n_233), .CI(n_56), .CO(n_61), .S(n_60));
   FA_X1 i_226 (.A(n_54), .B(n_43), .CI(n_41), .CO(n_63), .S(n_62));
   FA_X1 i_227 (.A(n_45), .B(n_60), .CI(n_58), .CO(n_65), .S(n_64));
   FA_X1 i_228 (.A(n_47), .B(n_62), .CI(n_49), .CO(n_67), .S(n_66));
   FA_X1 i_229 (.A(n_51), .B(n_64), .CI(n_66), .CO(n_69), .S(n_68));
   FA_X1 i_230 (.A(n_232), .B(n_231), .CI(n_230), .CO(n_71), .S(n_70));
   FA_X1 i_231 (.A(n_229), .B(n_55), .CI(n_228), .CO(n_73), .S(n_72));
   FA_X1 i_232 (.A(n_227), .B(n_226), .CI(n_225), .CO(n_75), .S(n_74));
   FA_X1 i_233 (.A(n_57), .B(n_70), .CI(n_59), .CO(n_77), .S(n_76));
   FA_X1 i_234 (.A(n_72), .B(n_63), .CI(n_61), .CO(n_79), .S(n_78));
   FA_X1 i_235 (.A(n_74), .B(n_76), .CI(n_65), .CO(n_81), .S(n_80));
   FA_X1 i_236 (.A(n_78), .B(n_67), .CI(n_80), .CO(n_83), .S(n_82));
   FA_X1 i_237 (.A(n_224), .B(n_223), .CI(n_222), .CO(n_85), .S(n_84));
   FA_X1 i_238 (.A(n_71), .B(n_221), .CI(n_220), .CO(n_87), .S(n_86));
   FA_X1 i_239 (.A(n_219), .B(n_218), .CI(n_84), .CO(n_89), .S(n_88));
   FA_X1 i_240 (.A(n_75), .B(n_73), .CI(n_77), .CO(n_91), .S(n_90));
   FA_X1 i_241 (.A(n_88), .B(n_86), .CI(n_79), .CO(n_93), .S(n_92));
   FA_X1 i_242 (.A(n_90), .B(n_81), .CI(n_92), .CO(n_95), .S(n_94));
   FA_X1 i_243 (.A(b_mantissa[14]), .B(n_217), .CI(n_216), .CO(n_97), .S(n_96));
   FA_X1 i_244 (.A(n_215), .B(n_85), .CI(n_214), .CO(n_99), .S(n_98));
   FA_X1 i_245 (.A(n_213), .B(n_212), .CI(n_211), .CO(n_101), .S(n_100));
   FA_X1 i_246 (.A(n_96), .B(n_87), .CI(n_98), .CO(n_103), .S(n_102));
   FA_X1 i_247 (.A(n_89), .B(n_100), .CI(n_91), .CO(n_105), .S(n_104));
   FA_X1 i_248 (.A(n_102), .B(n_93), .CI(n_104), .CO(n_107), .S(n_106));
   FA_X1 i_249 (.A(n_97), .B(n_210), .CI(n_209), .CO(n_109), .S(n_108));
   FA_X1 i_250 (.A(n_208), .B(n_99), .CI(n_1761), .CO(n_111), .S(n_110));
   FA_X1 i_251 (.A(n_101), .B(n_108), .CI(n_110), .CO(n_113), .S(n_112));
   FA_X1 i_252 (.A(n_103), .B(n_105), .CI(n_112), .CO(n_115), .S(n_114));
   FA_X1 i_253 (.A(n_207), .B(n_206), .CI(n_205), .CO(n_117), .S(n_116));
   FA_X1 i_254 (.A(n_1763), .B(n_109), .CI(n_111), .CO(n_119), .S(n_118));
   FA_X1 i_255 (.A(n_116), .B(n_118), .CI(n_113), .CO(n_121), .S(n_120));
   FA_X1 i_256 (.A(b_mantissa[17]), .B(n_204), .CI(n_203), .CO(n_123), .S(n_122));
   FA_X1 i_257 (.A(n_202), .B(n_201), .CI(n_200), .CO(n_125), .S(n_124));
   FA_X1 i_258 (.A(n_1764), .B(n_122), .CI(n_117), .CO(n_127), .S(n_126));
   FA_X1 i_259 (.A(n_124), .B(n_119), .CI(n_126), .CO(n_129), .S(n_128));
   FA_X1 i_260 (.A(n_199), .B(n_198), .CI(n_123), .CO(n_131), .S(n_130));
   FA_X1 i_261 (.A(n_197), .B(n_196), .CI(n_130), .CO(n_133), .S(n_132));
   FA_X1 i_262 (.A(n_125), .B(n_127), .CI(n_132), .CO(n_135), .S(n_134));
   FA_X1 i_263 (.A(n_131), .B(n_133), .CI(n_1838), .CO(n_137), .S(n_136));
   FA_X1 i_264 (.A(b_mantissa[20]), .B(n_195), .CI(n_194), .CO(n_139), .S(n_138));
   FA_X1 i_265 (.A(n_193), .B(n_138), .CI(n_1839), .CO(n_141), .S(n_140));
   FA_X1 i_266 (.A(n_192), .B(n_191), .CI(n_139), .CO(n_143), .S(n_142));
   FA_X1 i_267 (.A(a_mantissa[22]), .B(b_mantissa[22]), .CI(n_190), .CO(n_145), 
      .S(n_144));
   FA_X1 i_268 (.A(n_538), .B(n_533), .CI(n_189), .CO(n_146), .S(o_mantissa[3]));
   FA_X1 i_269 (.A(n_543), .B(n_556), .CI(n_146), .CO(n_147), .S(o_mantissa[4]));
   FA_X1 i_270 (.A(n_574), .B(n_572), .CI(n_147), .CO(n_148), .S(o_mantissa[5]));
   FA_X1 i_271 (.A(n_600), .B(n_598), .CI(n_148), .CO(n_149), .S(o_mantissa[6]));
   FA_X1 i_272 (.A(n_626), .B(n_628), .CI(n_149), .CO(n_150), .S(o_mantissa[7]));
   FA_X1 i_273 (.A(n_655), .B(n_657), .CI(n_150), .CO(n_151), .S(o_mantissa[8]));
   FA_X1 i_274 (.A(n_694), .B(n_692), .CI(n_151), .CO(n_152), .S(o_mantissa[9]));
   FA_X1 i_275 (.A(n_733), .B(n_731), .CI(n_152), .CO(n_153), .S(o_mantissa[10]));
   FA_X1 i_276 (.A(n_771), .B(n_773), .CI(n_153), .CO(n_154), .S(o_mantissa[11]));
   FA_X1 i_277 (.A(n_819), .B(n_821), .CI(n_154), .CO(n_155), .S(o_mantissa[12]));
   FA_X1 i_278 (.A(n_869), .B(n_871), .CI(n_155), .CO(n_156), .S(o_mantissa[13]));
   FA_X1 i_279 (.A(n_920), .B(n_922), .CI(n_156), .CO(n_157), .S(o_mantissa[14]));
   FA_X1 i_280 (.A(n_979), .B(n_981), .CI(n_157), .CO(n_158), .S(o_mantissa[15]));
   FA_X1 i_281 (.A(n_1040), .B(n_1042), .CI(n_158), .CO(n_159), .S(
      o_mantissa[16]));
   FA_X1 i_282 (.A(n_1102), .B(n_1104), .CI(n_159), .CO(n_160), .S(
      o_mantissa[17]));
   FA_X1 i_283 (.A(n_1105), .B(n_1174), .CI(n_160), .CO(n_161), .S(
      o_mantissa[18]));
   FA_X1 i_284 (.A(n_1175), .B(n_1246), .CI(n_161), .CO(n_162), .S(
      o_mantissa[19]));
   FA_X1 i_285 (.A(n_1317), .B(n_1319), .CI(n_162), .CO(n_163), .S(
      o_mantissa[20]));
   FA_X1 i_286 (.A(n_1320), .B(n_1400), .CI(n_163), .CO(n_164), .S(
      o_mantissa[21]));
   FA_X1 i_287 (.A(n_1401), .B(n_1483), .CI(n_164), .CO(n_165), .S(
      o_mantissa[22]));
   FA_X1 i_288 (.A(n_1484), .B(n_1569), .CI(n_165), .CO(n_166), .S(
      o_mantissa[23]));
   FA_X1 i_289 (.A(n_1570), .B(n_1655), .CI(n_166), .CO(n_167), .S(
      o_mantissa[24]));
   FA_X1 i_290 (.A(n_1656), .B(n_1733), .CI(n_167), .CO(n_168), .S(
      o_mantissa[25]));
   FA_X1 i_291 (.A(n_1734), .B(n_1810), .CI(n_168), .CO(n_169), .S(
      o_mantissa[26]));
   FA_X1 i_292 (.A(n_1811), .B(n_1885), .CI(n_169), .CO(n_170), .S(
      o_mantissa[27]));
   FA_X1 i_293 (.A(n_1886), .B(n_1952), .CI(n_170), .CO(n_171), .S(
      o_mantissa[28]));
   FA_X1 i_294 (.A(n_1953), .B(n_2018), .CI(n_171), .CO(n_172), .S(
      o_mantissa[29]));
   FA_X1 i_295 (.A(n_2019), .B(n_2082), .CI(n_172), .CO(n_173), .S(
      o_mantissa[30]));
   FA_X1 i_296 (.A(n_2083), .B(n_18), .CI(n_173), .CO(n_174), .S(o_mantissa[31]));
   FA_X1 i_297 (.A(n_19), .B(n_36), .CI(n_174), .CO(n_175), .S(o_mantissa[32]));
   FA_X1 i_298 (.A(n_52), .B(n_37), .CI(n_175), .CO(n_176), .S(o_mantissa[33]));
   FA_X1 i_299 (.A(n_53), .B(n_68), .CI(n_176), .CO(n_177), .S(o_mantissa[34]));
   FA_X1 i_300 (.A(n_69), .B(n_82), .CI(n_177), .CO(n_178), .S(o_mantissa[35]));
   FA_X1 i_301 (.A(n_94), .B(n_83), .CI(n_178), .CO(n_179), .S(o_mantissa[36]));
   FA_X1 i_302 (.A(n_95), .B(n_106), .CI(n_179), .CO(n_180), .S(o_mantissa[37]));
   FA_X1 i_303 (.A(n_107), .B(n_114), .CI(n_180), .CO(n_181), .S(o_mantissa[38]));
   FA_X1 i_304 (.A(n_120), .B(n_115), .CI(n_181), .CO(n_182), .S(o_mantissa[39]));
   FA_X1 i_305 (.A(n_121), .B(n_128), .CI(n_182), .CO(n_183), .S(o_mantissa[40]));
   FA_X1 i_306 (.A(n_134), .B(n_129), .CI(n_183), .CO(n_184), .S(o_mantissa[41]));
   FA_X1 i_307 (.A(n_135), .B(n_136), .CI(n_184), .CO(n_185), .S(o_mantissa[42]));
   FA_X1 i_308 (.A(n_140), .B(n_137), .CI(n_185), .CO(n_186), .S(o_mantissa[43]));
   FA_X1 i_309 (.A(n_141), .B(n_142), .CI(n_186), .CO(n_187), .S(o_mantissa[44]));
   FA_X1 i_310 (.A(n_144), .B(n_143), .CI(n_187), .CO(n_188), .S(o_mantissa[45]));
   XOR2_X1 i_311 (.A(n_2034), .B(n_248), .Z(n_543));
   NAND2_X1 i_312 (.A1(n_2039), .A2(n_2035), .ZN(n_248));
   AND2_X1 i_313 (.A1(n_2062), .A2(n_2057), .ZN(n_189));
   XOR2_X1 i_314 (.A(n_2053), .B(n_2049), .Z(n_533));
   XNOR2_X1 i_315 (.A(n_2089), .B(n_2048), .ZN(n_538));
   AOI22_X1 i_316 (.A1(n_1414), .A2(n_2111), .B1(n_1938), .B2(n_249), .ZN(n_190));
   XNOR2_X1 i_317 (.A(n_250), .B(n_249), .ZN(n_191));
   NAND2_X1 i_318 (.A1(b_mantissa[22]), .A2(a_mantissa[22]), .ZN(n_249));
   AOI21_X1 i_319 (.A(n_1901), .B1(n_1414), .B2(n_2111), .ZN(n_250));
   AOI21_X1 i_320 (.A(n_254), .B1(n_253), .B2(n_251), .ZN(n_192));
   XNOR2_X1 i_321 (.A(n_252), .B(n_251), .ZN(n_193));
   NAND2_X1 i_322 (.A1(b_mantissa[22]), .A2(a_mantissa[21]), .ZN(n_251));
   AOI21_X1 i_323 (.A(n_254), .B1(a_mantissa[22]), .B2(n_2107), .ZN(n_252));
   NAND2_X1 i_324 (.A1(a_mantissa[22]), .A2(n_2107), .ZN(n_253));
   AOI21_X1 i_325 (.A(a_mantissa[20]), .B1(b_mantissa[21]), .B2(a_mantissa[22]), 
      .ZN(n_254));
   AOI21_X1 i_326 (.A(n_2001), .B1(n_2008), .B2(n_1999), .ZN(n_194));
   AOI22_X1 i_327 (.A1(n_1198), .A2(n_1938), .B1(n_257), .B2(n_1900), .ZN(n_195));
   NAND2_X1 i_328 (.A1(a_mantissa[19]), .A2(n_1901), .ZN(n_257));
   XNOR2_X1 i_329 (.A(n_267), .B(n_2105), .ZN(n_196));
   AOI22_X1 i_330 (.A1(a_mantissa[18]), .A2(n_2107), .B1(n_1448), .B2(n_2110), 
      .ZN(n_267));
   XOR2_X1 i_331 (.A(n_273), .B(n_2098), .Z(n_197));
   OAI21_X1 i_332 (.A(n_2103), .B1(n_1409), .B2(n_2099), .ZN(n_273));
   AOI21_X1 i_333 (.A(n_280), .B1(n_278), .B2(n_276), .ZN(n_198));
   AOI22_X1 i_334 (.A1(n_294), .A2(n_2099), .B1(n_283), .B2(n_281), .ZN(n_199));
   XOR2_X1 i_335 (.A(n_277), .B(n_276), .Z(n_200));
   NAND2_X1 i_336 (.A1(b_mantissa[22]), .A2(a_mantissa[18]), .ZN(n_276));
   NAND2_X1 i_337 (.A1(n_279), .A2(n_278), .ZN(n_277));
   NAND3_X1 i_338 (.A1(b_mantissa[21]), .A2(a_mantissa[19]), .A3(a_mantissa[17]), 
      .ZN(n_278));
   INV_X1 i_339 (.A(n_280), .ZN(n_279));
   AOI21_X1 i_340 (.A(a_mantissa[17]), .B1(b_mantissa[21]), .B2(a_mantissa[19]), 
      .ZN(n_280));
   XNOR2_X1 i_341 (.A(n_282), .B(n_281), .ZN(n_201));
   NAND2_X1 i_342 (.A1(b_mantissa[20]), .A2(a_mantissa[20]), .ZN(n_281));
   AOI21_X1 i_343 (.A(n_284), .B1(n_294), .B2(n_2099), .ZN(n_282));
   INV_X1 i_344 (.A(n_284), .ZN(n_283));
   NOR2_X1 i_345 (.A1(n_294), .A2(n_2099), .ZN(n_284));
   AOI21_X1 i_346 (.A(n_299), .B1(n_300), .B2(n_296), .ZN(n_202));
   AOI21_X1 i_347 (.A(n_290), .B1(n_288), .B2(n_286), .ZN(n_203));
   OAI22_X1 i_348 (.A1(n_1835), .A2(n_294), .B1(n_295), .B2(n_291), .ZN(n_204));
   XOR2_X1 i_349 (.A(n_287), .B(n_286), .Z(n_205));
   NAND2_X1 i_350 (.A1(b_mantissa[22]), .A2(a_mantissa[17]), .ZN(n_286));
   NAND2_X1 i_351 (.A1(n_289), .A2(n_288), .ZN(n_287));
   NAND3_X1 i_352 (.A1(b_mantissa[21]), .A2(a_mantissa[18]), .A3(a_mantissa[16]), 
      .ZN(n_288));
   INV_X1 i_353 (.A(n_290), .ZN(n_289));
   AOI21_X1 i_354 (.A(a_mantissa[16]), .B1(b_mantissa[21]), .B2(a_mantissa[18]), 
      .ZN(n_290));
   XNOR2_X1 i_355 (.A(n_292), .B(n_291), .ZN(n_206));
   NAND2_X1 i_356 (.A1(b_mantissa[20]), .A2(a_mantissa[19]), .ZN(n_291));
   NOR2_X1 i_357 (.A1(n_295), .A2(n_293), .ZN(n_292));
   NOR2_X1 i_358 (.A1(n_1835), .A2(n_294), .ZN(n_293));
   NAND2_X1 i_359 (.A1(b_mantissa[19]), .A2(a_mantissa[21]), .ZN(n_294));
   AOI22_X1 i_360 (.A1(b_mantissa[19]), .A2(a_mantissa[20]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[21]), .ZN(n_295));
   XOR2_X1 i_361 (.A(n_297), .B(n_296), .Z(n_207));
   NAND2_X1 i_362 (.A1(b_mantissa[17]), .A2(a_mantissa[22]), .ZN(n_296));
   NAND2_X1 i_363 (.A1(n_300), .A2(n_298), .ZN(n_297));
   INV_X1 i_364 (.A(n_299), .ZN(n_298));
   AOI21_X1 i_365 (.A(b_mantissa[16]), .B1(b_mantissa[15]), .B2(n_313), .ZN(
      n_299));
   NAND2_X1 i_366 (.A1(n_316), .A2(n_301), .ZN(n_300));
   AOI21_X1 i_367 (.A(n_266), .B1(n_1816), .B2(n_314), .ZN(n_301));
   XOR2_X1 i_368 (.A(n_303), .B(n_1819), .Z(n_208));
   NAND2_X1 i_369 (.A1(n_305), .A2(n_1821), .ZN(n_303));
   INV_X1 i_370 (.A(n_1824), .ZN(n_305));
   XOR2_X1 i_371 (.A(n_308), .B(n_1827), .Z(n_209));
   NAND2_X1 i_372 (.A1(n_1831), .A2(n_1832), .ZN(n_308));
   XOR2_X1 i_373 (.A(n_315), .B(n_314), .Z(n_210));
   INV_X1 i_374 (.A(n_314), .ZN(n_313));
   NAND2_X1 i_375 (.A1(b_mantissa[17]), .A2(a_mantissa[21]), .ZN(n_314));
   OAI21_X1 i_376 (.A(n_316), .B1(n_266), .B2(n_1816), .ZN(n_315));
   INV_X1 i_377 (.A(n_317), .ZN(n_316));
   AOI21_X1 i_378 (.A(b_mantissa[15]), .B1(b_mantissa[16]), .B2(a_mantissa[22]), 
      .ZN(n_317));
   XNOR2_X1 i_379 (.A(n_319), .B(n_1765), .ZN(n_211));
   AOI21_X1 i_380 (.A(n_1768), .B1(a_mantissa[16]), .B2(n_357), .ZN(n_319));
   XOR2_X1 i_381 (.A(n_322), .B(n_1772), .Z(n_212));
   NAND2_X1 i_382 (.A1(n_324), .A2(n_1785), .ZN(n_322));
   INV_X1 i_383 (.A(n_1784), .ZN(n_324));
   XNOR2_X1 i_384 (.A(n_328), .B(n_1791), .ZN(n_213));
   AOI21_X1 i_385 (.A(n_1801), .B1(n_1818), .B2(n_1816), .ZN(n_328));
   AOI21_X1 i_386 (.A(n_351), .B1(n_352), .B2(n_348), .ZN(n_214));
   AOI21_X1 i_387 (.A(n_336), .B1(n_334), .B2(n_332), .ZN(n_215));
   OAI21_X1 i_388 (.A(n_339), .B1(n_340), .B2(n_337), .ZN(n_216));
   OAI22_X1 i_389 (.A1(n_370), .A2(n_1818), .B1(n_347), .B2(n_343), .ZN(n_217));
   XOR2_X1 i_390 (.A(n_333), .B(n_332), .Z(n_218));
   NAND2_X1 i_391 (.A1(b_mantissa[22]), .A2(a_mantissa[14]), .ZN(n_332));
   NAND2_X1 i_392 (.A1(n_335), .A2(n_334), .ZN(n_333));
   NAND3_X1 i_393 (.A1(b_mantissa[21]), .A2(a_mantissa[15]), .A3(a_mantissa[13]), 
      .ZN(n_334));
   INV_X1 i_394 (.A(n_336), .ZN(n_335));
   AOI21_X1 i_395 (.A(a_mantissa[13]), .B1(b_mantissa[21]), .B2(a_mantissa[15]), 
      .ZN(n_336));
   XOR2_X1 i_396 (.A(n_338), .B(n_337), .Z(n_219));
   NAND2_X1 i_397 (.A1(b_mantissa[20]), .A2(a_mantissa[16]), .ZN(n_337));
   NAND2_X1 i_398 (.A1(n_341), .A2(n_339), .ZN(n_338));
   OR3_X1 i_399 (.A1(n_1409), .A2(n_2106), .A3(n_342), .ZN(n_339));
   INV_X1 i_400 (.A(n_341), .ZN(n_340));
   OAI21_X1 i_401 (.A(n_342), .B1(n_1409), .B2(n_2106), .ZN(n_341));
   NAND2_X1 i_402 (.A1(b_mantissa[18]), .A2(a_mantissa[18]), .ZN(n_342));
   XNOR2_X1 i_403 (.A(n_344), .B(n_343), .ZN(n_220));
   NAND2_X1 i_404 (.A1(b_mantissa[17]), .A2(a_mantissa[19]), .ZN(n_343));
   NOR2_X1 i_405 (.A1(n_347), .A2(n_345), .ZN(n_344));
   NOR2_X1 i_406 (.A1(n_370), .A2(n_1818), .ZN(n_345));
   AOI22_X1 i_407 (.A1(b_mantissa[16]), .A2(a_mantissa[20]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[21]), .ZN(n_347));
   XOR2_X1 i_408 (.A(n_349), .B(n_348), .Z(n_221));
   NAND2_X1 i_409 (.A1(b_mantissa[14]), .A2(a_mantissa[22]), .ZN(n_348));
   NAND2_X1 i_410 (.A1(n_352), .A2(n_350), .ZN(n_349));
   INV_X1 i_411 (.A(n_351), .ZN(n_350));
   AOI21_X1 i_412 (.A(b_mantissa[13]), .B1(b_mantissa[12]), .B2(n_371), .ZN(
      n_351));
   NAND2_X1 i_413 (.A1(n_374), .A2(n_353), .ZN(n_352));
   AOI21_X1 i_414 (.A(n_1506), .B1(n_396), .B2(n_372), .ZN(n_353));
   AOI22_X1 i_415 (.A1(n_1507), .A2(n_1770), .B1(n_356), .B2(n_354), .ZN(n_222));
   OAI21_X1 i_416 (.A(n_361), .B1(n_362), .B2(n_359), .ZN(n_223));
   OAI21_X1 i_417 (.A(n_367), .B1(n_368), .B2(n_365), .ZN(n_224));
   XNOR2_X1 i_418 (.A(n_355), .B(n_354), .ZN(n_225));
   NAND2_X1 i_419 (.A1(b_mantissa[22]), .A2(a_mantissa[13]), .ZN(n_354));
   AOI22_X1 i_420 (.A1(a_mantissa[12]), .A2(n_357), .B1(n_1507), .B2(n_1770), 
      .ZN(n_355));
   NAND2_X1 i_421 (.A1(a_mantissa[12]), .A2(n_357), .ZN(n_356));
   INV_X1 i_422 (.A(n_1770), .ZN(n_357));
   XOR2_X1 i_423 (.A(n_360), .B(n_359), .Z(n_226));
   NAND2_X1 i_424 (.A1(b_mantissa[20]), .A2(a_mantissa[15]), .ZN(n_359));
   NAND2_X1 i_425 (.A1(n_363), .A2(n_361), .ZN(n_360));
   OR3_X1 i_426 (.A1(n_1409), .A2(n_957), .A3(n_364), .ZN(n_361));
   INV_X1 i_427 (.A(n_363), .ZN(n_362));
   OAI21_X1 i_428 (.A(n_364), .B1(n_1409), .B2(n_957), .ZN(n_363));
   NAND2_X1 i_429 (.A1(b_mantissa[18]), .A2(a_mantissa[17]), .ZN(n_364));
   XOR2_X1 i_430 (.A(n_366), .B(n_365), .Z(n_227));
   NAND2_X1 i_431 (.A1(b_mantissa[17]), .A2(a_mantissa[18]), .ZN(n_365));
   NAND2_X1 i_432 (.A1(n_369), .A2(n_367), .ZN(n_366));
   NAND3_X1 i_433 (.A1(b_mantissa[16]), .A2(a_mantissa[20]), .A3(n_391), 
      .ZN(n_367));
   INV_X1 i_434 (.A(n_369), .ZN(n_368));
   OAI21_X1 i_435 (.A(n_370), .B1(n_266), .B2(n_1198), .ZN(n_369));
   NAND2_X1 i_436 (.A1(b_mantissa[15]), .A2(a_mantissa[20]), .ZN(n_370));
   XOR2_X1 i_437 (.A(n_373), .B(n_372), .Z(n_228));
   INV_X1 i_438 (.A(n_372), .ZN(n_371));
   NAND2_X1 i_439 (.A1(b_mantissa[14]), .A2(a_mantissa[21]), .ZN(n_372));
   OAI21_X1 i_440 (.A(n_374), .B1(n_1506), .B2(n_396), .ZN(n_373));
   INV_X1 i_441 (.A(n_375), .ZN(n_374));
   AOI21_X1 i_442 (.A(b_mantissa[12]), .B1(b_mantissa[13]), .B2(a_mantissa[22]), 
      .ZN(n_375));
   AOI21_X1 i_443 (.A(n_380), .B1(n_378), .B2(n_376), .ZN(n_229));
   OAI21_X1 i_444 (.A(n_383), .B1(n_385), .B2(n_381), .ZN(n_230));
   OAI21_X1 i_445 (.A(n_388), .B1(n_390), .B2(n_386), .ZN(n_231));
   OAI22_X1 i_446 (.A1(n_416), .A2(n_396), .B1(n_394), .B2(n_392), .ZN(n_232));
   XOR2_X1 i_447 (.A(n_377), .B(n_376), .Z(n_233));
   NAND2_X1 i_448 (.A1(b_mantissa[22]), .A2(a_mantissa[12]), .ZN(n_376));
   NAND2_X1 i_449 (.A1(n_379), .A2(n_378), .ZN(n_377));
   NAND3_X1 i_450 (.A1(b_mantissa[21]), .A2(a_mantissa[13]), .A3(a_mantissa[11]), 
      .ZN(n_378));
   INV_X1 i_451 (.A(n_380), .ZN(n_379));
   AOI21_X1 i_452 (.A(a_mantissa[11]), .B1(b_mantissa[21]), .B2(a_mantissa[13]), 
      .ZN(n_380));
   XOR2_X1 i_453 (.A(n_382), .B(n_381), .Z(n_234));
   NAND2_X1 i_454 (.A1(b_mantissa[20]), .A2(a_mantissa[14]), .ZN(n_381));
   NAND2_X1 i_455 (.A1(n_384), .A2(n_383), .ZN(n_382));
   NAND3_X1 i_456 (.A1(b_mantissa[18]), .A2(a_mantissa[16]), .A3(n_405), 
      .ZN(n_383));
   INV_X1 i_457 (.A(n_385), .ZN(n_384));
   AOI21_X1 i_458 (.A(n_405), .B1(b_mantissa[18]), .B2(a_mantissa[16]), .ZN(
      n_385));
   XOR2_X1 i_459 (.A(n_387), .B(n_386), .Z(n_235));
   NAND2_X1 i_460 (.A1(b_mantissa[17]), .A2(a_mantissa[17]), .ZN(n_386));
   NAND2_X1 i_461 (.A1(n_389), .A2(n_388), .ZN(n_387));
   NAND3_X1 i_462 (.A1(b_mantissa[16]), .A2(a_mantissa[18]), .A3(n_391), 
      .ZN(n_388));
   INV_X1 i_463 (.A(n_390), .ZN(n_389));
   AOI21_X1 i_464 (.A(n_391), .B1(b_mantissa[16]), .B2(a_mantissa[18]), .ZN(
      n_390));
   AND2_X1 i_465 (.A1(b_mantissa[15]), .A2(a_mantissa[19]), .ZN(n_391));
   XOR2_X1 i_466 (.A(n_393), .B(n_392), .Z(n_236));
   NAND2_X1 i_467 (.A1(b_mantissa[14]), .A2(a_mantissa[20]), .ZN(n_392));
   OAI21_X1 i_468 (.A(n_395), .B1(n_416), .B2(n_396), .ZN(n_393));
   INV_X1 i_469 (.A(n_395), .ZN(n_394));
   NAND2_X1 i_470 (.A1(n_416), .A2(n_396), .ZN(n_395));
   NAND2_X1 i_471 (.A1(b_mantissa[12]), .A2(a_mantissa[22]), .ZN(n_396));
   AOI21_X1 i_472 (.A(n_422), .B1(n_423), .B2(n_419), .ZN(n_237));
   AOI21_X1 i_473 (.A(n_401), .B1(n_399), .B2(n_397), .ZN(n_238));
   OAI21_X1 i_474 (.A(n_404), .B1(n_407), .B2(n_402), .ZN(n_239));
   OAI21_X1 i_475 (.A(n_410), .B1(n_411), .B2(n_408), .ZN(n_240));
   OAI22_X1 i_476 (.A1(n_446), .A2(n_416), .B1(n_418), .B2(n_414), .ZN(n_241));
   XOR2_X1 i_477 (.A(n_398), .B(n_397), .Z(n_242));
   NAND2_X1 i_478 (.A1(b_mantissa[22]), .A2(a_mantissa[11]), .ZN(n_397));
   NAND2_X1 i_479 (.A1(n_400), .A2(n_399), .ZN(n_398));
   NAND3_X1 i_480 (.A1(b_mantissa[21]), .A2(a_mantissa[12]), .A3(a_mantissa[10]), 
      .ZN(n_399));
   INV_X1 i_481 (.A(n_401), .ZN(n_400));
   AOI21_X1 i_482 (.A(a_mantissa[10]), .B1(b_mantissa[21]), .B2(a_mantissa[12]), 
      .ZN(n_401));
   XOR2_X1 i_483 (.A(n_403), .B(n_402), .Z(n_243));
   NAND2_X1 i_484 (.A1(b_mantissa[20]), .A2(a_mantissa[13]), .ZN(n_402));
   NAND2_X1 i_485 (.A1(n_406), .A2(n_404), .ZN(n_403));
   NAND3_X1 i_486 (.A1(b_mantissa[18]), .A2(a_mantissa[14]), .A3(n_405), 
      .ZN(n_404));
   NOR2_X1 i_487 (.A1(n_1409), .A2(n_1518), .ZN(n_405));
   INV_X1 i_488 (.A(n_407), .ZN(n_406));
   AOI22_X1 i_489 (.A1(b_mantissa[19]), .A2(a_mantissa[14]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[15]), .ZN(n_407));
   XOR2_X1 i_490 (.A(n_409), .B(n_408), .Z(n_244));
   NAND2_X1 i_491 (.A1(b_mantissa[17]), .A2(a_mantissa[16]), .ZN(n_408));
   NAND2_X1 i_492 (.A1(n_412), .A2(n_410), .ZN(n_409));
   OR3_X1 i_493 (.A1(n_266), .A2(n_2106), .A3(n_413), .ZN(n_410));
   INV_X1 i_494 (.A(n_412), .ZN(n_411));
   OAI21_X1 i_495 (.A(n_413), .B1(n_266), .B2(n_2106), .ZN(n_412));
   NAND2_X1 i_496 (.A1(b_mantissa[15]), .A2(a_mantissa[18]), .ZN(n_413));
   XOR2_X1 i_497 (.A(n_415), .B(n_414), .Z(n_245));
   NAND2_X1 i_498 (.A1(b_mantissa[14]), .A2(a_mantissa[19]), .ZN(n_414));
   OAI21_X1 i_499 (.A(n_417), .B1(n_446), .B2(n_416), .ZN(n_415));
   NAND2_X1 i_500 (.A1(b_mantissa[13]), .A2(a_mantissa[21]), .ZN(n_416));
   INV_X1 i_501 (.A(n_418), .ZN(n_417));
   AOI22_X1 i_502 (.A1(b_mantissa[13]), .A2(a_mantissa[20]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[21]), .ZN(n_418));
   XOR2_X1 i_503 (.A(n_420), .B(n_419), .Z(n_246));
   NAND2_X1 i_504 (.A1(b_mantissa[11]), .A2(a_mantissa[22]), .ZN(n_419));
   NAND2_X1 i_505 (.A1(n_423), .A2(n_421), .ZN(n_420));
   INV_X1 i_506 (.A(n_422), .ZN(n_421));
   AOI21_X1 i_507 (.A(b_mantissa[10]), .B1(b_mantissa[9]), .B2(n_447), .ZN(n_422));
   NAND2_X1 i_508 (.A1(n_450), .A2(n_424), .ZN(n_423));
   AOI21_X1 i_509 (.A(n_554), .B1(n_476), .B2(n_448), .ZN(n_424));
   AOI21_X1 i_510 (.A(n_429), .B1(n_427), .B2(n_425), .ZN(n_247));
   OAI21_X1 i_511 (.A(n_432), .B1(n_434), .B2(n_430), .ZN(n_255));
   OAI21_X1 i_512 (.A(n_437), .B1(n_438), .B2(n_435), .ZN(n_256));
   OAI21_X1 i_513 (.A(n_443), .B1(n_444), .B2(n_441), .ZN(n_258));
   XOR2_X1 i_514 (.A(n_426), .B(n_425), .Z(n_259));
   NAND2_X1 i_515 (.A1(b_mantissa[22]), .A2(a_mantissa[10]), .ZN(n_425));
   NAND2_X1 i_516 (.A1(n_428), .A2(n_427), .ZN(n_426));
   NAND3_X1 i_517 (.A1(b_mantissa[21]), .A2(a_mantissa[11]), .A3(a_mantissa[9]), 
      .ZN(n_427));
   INV_X1 i_518 (.A(n_429), .ZN(n_428));
   AOI21_X1 i_519 (.A(a_mantissa[9]), .B1(b_mantissa[21]), .B2(a_mantissa[11]), 
      .ZN(n_429));
   XOR2_X1 i_520 (.A(n_431), .B(n_430), .Z(n_260));
   NAND2_X1 i_521 (.A1(b_mantissa[20]), .A2(a_mantissa[12]), .ZN(n_430));
   NAND2_X1 i_522 (.A1(n_433), .A2(n_432), .ZN(n_431));
   NAND4_X1 i_523 (.A1(b_mantissa[18]), .A2(a_mantissa[13]), .A3(b_mantissa[19]), 
      .A4(a_mantissa[14]), .ZN(n_432));
   INV_X1 i_524 (.A(n_434), .ZN(n_433));
   AOI22_X1 i_525 (.A1(b_mantissa[19]), .A2(a_mantissa[13]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[14]), .ZN(n_434));
   XOR2_X1 i_526 (.A(n_436), .B(n_435), .Z(n_261));
   NAND2_X1 i_527 (.A1(b_mantissa[17]), .A2(a_mantissa[15]), .ZN(n_435));
   NAND2_X1 i_528 (.A1(n_439), .A2(n_437), .ZN(n_436));
   OR3_X1 i_529 (.A1(n_266), .A2(n_957), .A3(n_440), .ZN(n_437));
   INV_X1 i_530 (.A(n_439), .ZN(n_438));
   OAI21_X1 i_531 (.A(n_440), .B1(n_266), .B2(n_957), .ZN(n_439));
   NAND2_X1 i_532 (.A1(b_mantissa[15]), .A2(a_mantissa[17]), .ZN(n_440));
   XOR2_X1 i_533 (.A(n_442), .B(n_441), .Z(n_262));
   NAND2_X1 i_534 (.A1(b_mantissa[14]), .A2(a_mantissa[18]), .ZN(n_441));
   NAND2_X1 i_535 (.A1(n_445), .A2(n_443), .ZN(n_442));
   OR3_X1 i_536 (.A1(n_1506), .A2(n_1198), .A3(n_446), .ZN(n_443));
   INV_X1 i_537 (.A(n_445), .ZN(n_444));
   OAI21_X1 i_538 (.A(n_446), .B1(n_1506), .B2(n_1198), .ZN(n_445));
   NAND2_X1 i_539 (.A1(b_mantissa[12]), .A2(a_mantissa[20]), .ZN(n_446));
   XOR2_X1 i_540 (.A(n_449), .B(n_448), .Z(n_263));
   INV_X1 i_541 (.A(n_448), .ZN(n_447));
   NAND2_X1 i_542 (.A1(b_mantissa[11]), .A2(a_mantissa[21]), .ZN(n_448));
   OAI21_X1 i_543 (.A(n_450), .B1(n_554), .B2(n_476), .ZN(n_449));
   INV_X1 i_544 (.A(n_451), .ZN(n_450));
   AOI21_X1 i_545 (.A(b_mantissa[9]), .B1(b_mantissa[10]), .B2(a_mantissa[22]), 
      .ZN(n_451));
   AOI21_X1 i_546 (.A(n_456), .B1(n_454), .B2(n_452), .ZN(n_2086));
   AOI22_X1 i_547 (.A1(n_484), .A2(n_461), .B1(n_460), .B2(n_457), .ZN(n_2095));
   OAI21_X1 i_548 (.A(n_464), .B1(n_466), .B2(n_462), .ZN(n_2102));
   OAI22_X1 i_549 (.A1(n_495), .A2(n_471), .B1(n_469), .B2(n_467), .ZN(n_2109));
   AOI22_X1 i_550 (.A1(n_501), .A2(n_476), .B1(n_474), .B2(n_472), .ZN(n_264));
   XOR2_X1 i_551 (.A(n_453), .B(n_452), .Z(n_2085));
   NAND2_X1 i_552 (.A1(b_mantissa[22]), .A2(a_mantissa[9]), .ZN(n_452));
   NAND2_X1 i_553 (.A1(n_455), .A2(n_454), .ZN(n_453));
   NAND3_X1 i_554 (.A1(b_mantissa[21]), .A2(a_mantissa[10]), .A3(a_mantissa[8]), 
      .ZN(n_454));
   INV_X1 i_555 (.A(n_456), .ZN(n_455));
   AOI21_X1 i_556 (.A(a_mantissa[8]), .B1(b_mantissa[21]), .B2(a_mantissa[10]), 
      .ZN(n_456));
   XOR2_X1 i_557 (.A(n_458), .B(n_457), .Z(n_2094));
   NAND2_X1 i_558 (.A1(b_mantissa[20]), .A2(a_mantissa[11]), .ZN(n_457));
   NAND2_X1 i_559 (.A1(n_460), .A2(n_459), .ZN(n_458));
   NAND2_X1 i_560 (.A1(n_484), .A2(n_461), .ZN(n_459));
   OR2_X1 i_561 (.A1(n_484), .A2(n_461), .ZN(n_460));
   NAND2_X1 i_562 (.A1(b_mantissa[18]), .A2(a_mantissa[13]), .ZN(n_461));
   XOR2_X1 i_563 (.A(n_463), .B(n_462), .Z(n_2101));
   NAND2_X1 i_564 (.A1(b_mantissa[17]), .A2(a_mantissa[14]), .ZN(n_462));
   NAND2_X1 i_565 (.A1(n_465), .A2(n_464), .ZN(n_463));
   NAND3_X1 i_566 (.A1(b_mantissa[15]), .A2(a_mantissa[16]), .A3(n_490), 
      .ZN(n_464));
   INV_X1 i_567 (.A(n_466), .ZN(n_465));
   AOI21_X1 i_568 (.A(n_490), .B1(b_mantissa[15]), .B2(a_mantissa[16]), .ZN(
      n_466));
   XOR2_X1 i_569 (.A(n_468), .B(n_467), .Z(n_2108));
   NAND2_X1 i_570 (.A1(b_mantissa[14]), .A2(a_mantissa[17]), .ZN(n_467));
   OAI21_X1 i_571 (.A(n_470), .B1(n_495), .B2(n_471), .ZN(n_468));
   INV_X1 i_572 (.A(n_470), .ZN(n_469));
   NAND2_X1 i_573 (.A1(n_495), .A2(n_471), .ZN(n_470));
   NAND2_X1 i_574 (.A1(b_mantissa[12]), .A2(a_mantissa[19]), .ZN(n_471));
   XNOR2_X1 i_575 (.A(n_473), .B(n_472), .ZN(n_265));
   NAND2_X1 i_576 (.A1(b_mantissa[11]), .A2(a_mantissa[20]), .ZN(n_472));
   AOI21_X1 i_577 (.A(n_475), .B1(n_501), .B2(n_476), .ZN(n_473));
   INV_X1 i_578 (.A(n_475), .ZN(n_474));
   NOR2_X1 i_579 (.A1(n_501), .A2(n_476), .ZN(n_475));
   NAND2_X1 i_580 (.A1(b_mantissa[9]), .A2(a_mantissa[22]), .ZN(n_476));
   AOI21_X1 i_581 (.A(n_506), .B1(n_507), .B2(n_503), .ZN(n_2059));
   AOI21_X1 i_582 (.A(n_481), .B1(n_479), .B2(n_477), .ZN(n_2022));
   OAI22_X1 i_583 (.A1(n_519), .A2(n_484), .B1(n_486), .B2(n_482), .ZN(n_2031));
   OAI21_X1 i_584 (.A(n_489), .B1(n_492), .B2(n_487), .ZN(n_2038));
   OAI22_X1 i_585 (.A1(n_530), .A2(n_495), .B1(n_497), .B2(n_493), .ZN(n_2045));
   OAI22_X1 i_586 (.A1(n_539), .A2(n_501), .B1(n_502), .B2(n_498), .ZN(n_2052));
   XOR2_X1 i_587 (.A(n_478), .B(n_477), .Z(n_2021));
   NAND2_X1 i_588 (.A1(b_mantissa[22]), .A2(a_mantissa[8]), .ZN(n_477));
   NAND2_X1 i_589 (.A1(n_480), .A2(n_479), .ZN(n_478));
   NAND3_X1 i_590 (.A1(b_mantissa[21]), .A2(a_mantissa[9]), .A3(a_mantissa[7]), 
      .ZN(n_479));
   INV_X1 i_591 (.A(n_481), .ZN(n_480));
   AOI21_X1 i_592 (.A(a_mantissa[7]), .B1(b_mantissa[21]), .B2(a_mantissa[9]), 
      .ZN(n_481));
   XOR2_X1 i_593 (.A(n_483), .B(n_482), .Z(n_2030));
   NAND2_X1 i_594 (.A1(b_mantissa[20]), .A2(a_mantissa[10]), .ZN(n_482));
   OAI21_X1 i_595 (.A(n_485), .B1(n_519), .B2(n_484), .ZN(n_483));
   NAND2_X1 i_596 (.A1(b_mantissa[19]), .A2(a_mantissa[12]), .ZN(n_484));
   INV_X1 i_597 (.A(n_486), .ZN(n_485));
   AOI22_X1 i_598 (.A1(b_mantissa[19]), .A2(a_mantissa[11]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[12]), .ZN(n_486));
   XOR2_X1 i_599 (.A(n_488), .B(n_487), .Z(n_2037));
   NAND2_X1 i_600 (.A1(b_mantissa[17]), .A2(a_mantissa[13]), .ZN(n_487));
   NAND2_X1 i_601 (.A1(n_491), .A2(n_489), .ZN(n_488));
   NAND3_X1 i_602 (.A1(b_mantissa[15]), .A2(a_mantissa[14]), .A3(n_490), 
      .ZN(n_489));
   NOR2_X1 i_603 (.A1(n_266), .A2(n_1518), .ZN(n_490));
   INV_X1 i_604 (.A(n_492), .ZN(n_491));
   AOI22_X1 i_605 (.A1(b_mantissa[16]), .A2(a_mantissa[14]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[15]), .ZN(n_492));
   XOR2_X1 i_606 (.A(n_494), .B(n_493), .Z(n_2044));
   NAND2_X1 i_607 (.A1(b_mantissa[14]), .A2(a_mantissa[16]), .ZN(n_493));
   OAI21_X1 i_608 (.A(n_496), .B1(n_530), .B2(n_495), .ZN(n_494));
   NAND2_X1 i_609 (.A1(b_mantissa[13]), .A2(a_mantissa[18]), .ZN(n_495));
   INV_X1 i_610 (.A(n_497), .ZN(n_496));
   AOI22_X1 i_611 (.A1(b_mantissa[13]), .A2(a_mantissa[17]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[18]), .ZN(n_497));
   XNOR2_X1 i_612 (.A(n_499), .B(n_498), .ZN(n_2051));
   NAND2_X1 i_613 (.A1(b_mantissa[11]), .A2(a_mantissa[19]), .ZN(n_498));
   NOR2_X1 i_614 (.A1(n_502), .A2(n_500), .ZN(n_499));
   NOR2_X1 i_615 (.A1(n_539), .A2(n_501), .ZN(n_500));
   NAND2_X1 i_616 (.A1(b_mantissa[10]), .A2(a_mantissa[21]), .ZN(n_501));
   AOI22_X1 i_617 (.A1(b_mantissa[10]), .A2(a_mantissa[20]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[21]), .ZN(n_502));
   XOR2_X1 i_618 (.A(n_504), .B(n_503), .Z(n_2058));
   NAND2_X1 i_619 (.A1(b_mantissa[8]), .A2(a_mantissa[22]), .ZN(n_503));
   NAND2_X1 i_620 (.A1(n_507), .A2(n_505), .ZN(n_504));
   INV_X1 i_621 (.A(n_506), .ZN(n_505));
   AOI21_X1 i_622 (.A(b_mantissa[7]), .B1(b_mantissa[6]), .B2(n_540), .ZN(n_506));
   OAI21_X1 i_623 (.A(n_508), .B1(n_1740), .B2(n_540), .ZN(n_507));
   NOR2_X1 i_624 (.A1(n_1445), .A2(n_542), .ZN(n_508));
   AOI21_X1 i_625 (.A(n_513), .B1(n_511), .B2(n_509), .ZN(n_1956));
   OAI21_X1 i_626 (.A(n_518), .B1(n_516), .B2(n_514), .ZN(n_1965));
   OAI21_X1 i_627 (.A(n_524), .B1(n_523), .B2(n_520), .ZN(n_1972));
   OAI21_X1 i_628 (.A(n_527), .B1(n_528), .B2(n_525), .ZN(n_1979));
   OAI21_X1 i_629 (.A(n_535), .B1(n_536), .B2(n_531), .ZN(n_1986));
   XOR2_X1 i_630 (.A(n_510), .B(n_509), .Z(n_1955));
   NAND2_X1 i_631 (.A1(b_mantissa[22]), .A2(a_mantissa[7]), .ZN(n_509));
   NAND2_X1 i_632 (.A1(n_512), .A2(n_511), .ZN(n_510));
   NAND3_X1 i_633 (.A1(b_mantissa[21]), .A2(a_mantissa[8]), .A3(a_mantissa[6]), 
      .ZN(n_511));
   INV_X1 i_634 (.A(n_513), .ZN(n_512));
   AOI21_X1 i_635 (.A(a_mantissa[6]), .B1(b_mantissa[21]), .B2(a_mantissa[8]), 
      .ZN(n_513));
   XOR2_X1 i_636 (.A(n_515), .B(n_514), .Z(n_1964));
   NAND2_X1 i_637 (.A1(b_mantissa[20]), .A2(a_mantissa[9]), .ZN(n_514));
   NAND2_X1 i_638 (.A1(n_518), .A2(n_517), .ZN(n_515));
   INV_X1 i_639 (.A(n_517), .ZN(n_516));
   OAI21_X1 i_640 (.A(n_519), .B1(n_1409), .B2(n_2100), .ZN(n_517));
   NAND3_X1 i_641 (.A1(b_mantissa[19]), .A2(a_mantissa[11]), .A3(n_1754), 
      .ZN(n_518));
   NAND2_X1 i_642 (.A1(b_mantissa[18]), .A2(a_mantissa[11]), .ZN(n_519));
   XOR2_X1 i_643 (.A(n_521), .B(n_520), .Z(n_1971));
   NAND2_X1 i_644 (.A1(b_mantissa[17]), .A2(a_mantissa[12]), .ZN(n_520));
   NAND2_X1 i_645 (.A1(n_524), .A2(n_522), .ZN(n_521));
   INV_X1 i_646 (.A(n_523), .ZN(n_522));
   AOI22_X1 i_647 (.A1(b_mantissa[16]), .A2(a_mantissa[13]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[14]), .ZN(n_523));
   NAND3_X1 i_648 (.A1(b_mantissa[16]), .A2(a_mantissa[14]), .A3(n_1756), 
      .ZN(n_524));
   XOR2_X1 i_649 (.A(n_526), .B(n_525), .Z(n_1978));
   NAND2_X1 i_650 (.A1(b_mantissa[14]), .A2(a_mantissa[15]), .ZN(n_525));
   NAND2_X1 i_651 (.A1(n_529), .A2(n_527), .ZN(n_526));
   NAND3_X1 i_652 (.A1(b_mantissa[13]), .A2(a_mantissa[17]), .A3(n_1691), 
      .ZN(n_527));
   INV_X1 i_653 (.A(n_529), .ZN(n_528));
   OAI21_X1 i_654 (.A(n_530), .B1(n_1506), .B2(n_957), .ZN(n_529));
   NAND2_X1 i_655 (.A1(b_mantissa[12]), .A2(a_mantissa[17]), .ZN(n_530));
   XOR2_X1 i_656 (.A(n_532), .B(n_531), .Z(n_1985));
   NAND2_X1 i_657 (.A1(b_mantissa[11]), .A2(a_mantissa[18]), .ZN(n_531));
   NAND2_X1 i_658 (.A1(n_537), .A2(n_535), .ZN(n_532));
   NAND3_X1 i_659 (.A1(b_mantissa[10]), .A2(a_mantissa[20]), .A3(n_1735), 
      .ZN(n_535));
   INV_X1 i_660 (.A(n_537), .ZN(n_536));
   OAI21_X1 i_661 (.A(n_539), .B1(n_554), .B2(n_1198), .ZN(n_537));
   NAND2_X1 i_662 (.A1(b_mantissa[9]), .A2(a_mantissa[20]), .ZN(n_539));
   XOR2_X1 i_663 (.A(n_541), .B(n_540), .Z(n_1991));
   AND2_X1 i_664 (.A1(b_mantissa[8]), .A2(a_mantissa[21]), .ZN(n_540));
   AOI21_X1 i_665 (.A(n_542), .B1(b_mantissa[7]), .B2(n_1740), .ZN(n_541));
   AOI21_X1 i_666 (.A(b_mantissa[6]), .B1(b_mantissa[7]), .B2(a_mantissa[22]), 
      .ZN(n_542));
   XOR2_X1 i_667 (.A(n_548), .B(n_1748), .Z(n_1888));
   NAND2_X1 i_668 (.A1(n_552), .A2(n_1750), .ZN(n_548));
   INV_X1 i_669 (.A(n_1751), .ZN(n_552));
   XOR2_X1 i_670 (.A(n_582), .B(n_1709), .Z(n_1918));
   NAND2_X1 i_671 (.A1(n_584), .A2(n_1721), .ZN(n_582));
   INV_X1 i_672 (.A(n_1713), .ZN(n_584));
   XNOR2_X1 i_673 (.A(n_589), .B(n_1738), .ZN(n_1925));
   AOI22_X1 i_674 (.A1(n_1743), .A2(n_1740), .B1(n_1744), .B2(n_1742), .ZN(n_589));
   AOI21_X1 i_675 (.A(n_666), .B1(n_667), .B2(n_663), .ZN(n_1858));
   AOI21_X1 i_676 (.A(n_1621), .B1(n_1620), .B2(n_1619), .ZN(n_1814));
   OAI21_X1 i_677 (.A(n_1627), .B1(n_1626), .B2(n_1625), .ZN(n_1823));
   OAI21_X1 i_678 (.A(n_1660), .B1(n_1657), .B2(n_1637), .ZN(n_1830));
   OAI21_X1 i_679 (.A(n_634), .B1(n_638), .B2(n_630), .ZN(n_1837));
   OAI21_X1 i_680 (.A(n_642), .B1(n_643), .B2(n_640), .ZN(n_1844));
   AOI21_X1 i_681 (.A(n_660), .B1(n_649), .B2(n_647), .ZN(n_1851));
   XOR2_X1 i_682 (.A(n_631), .B(n_630), .Z(n_1836));
   NAND2_X1 i_683 (.A1(b_mantissa[14]), .A2(a_mantissa[13]), .ZN(n_630));
   NAND2_X1 i_684 (.A1(n_637), .A2(n_634), .ZN(n_631));
   NAND2_X1 i_685 (.A1(n_707), .A2(n_1704), .ZN(n_634));
   INV_X1 i_686 (.A(n_638), .ZN(n_637));
   AOI22_X1 i_687 (.A1(b_mantissa[13]), .A2(a_mantissa[14]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[15]), .ZN(n_638));
   XOR2_X1 i_688 (.A(n_641), .B(n_640), .Z(n_1843));
   NAND2_X1 i_689 (.A1(b_mantissa[11]), .A2(a_mantissa[16]), .ZN(n_640));
   NAND2_X1 i_690 (.A1(n_644), .A2(n_642), .ZN(n_641));
   OR3_X1 i_691 (.A1(n_554), .A2(n_2106), .A3(n_645), .ZN(n_642));
   INV_X1 i_692 (.A(n_644), .ZN(n_643));
   OAI21_X1 i_693 (.A(n_645), .B1(n_554), .B2(n_2106), .ZN(n_644));
   NAND2_X1 i_694 (.A1(b_mantissa[9]), .A2(a_mantissa[18]), .ZN(n_645));
   XNOR2_X1 i_695 (.A(n_648), .B(n_647), .ZN(n_1850));
   NAND2_X1 i_696 (.A1(b_mantissa[8]), .A2(a_mantissa[19]), .ZN(n_647));
   AOI21_X1 i_697 (.A(n_660), .B1(n_723), .B2(n_1743), .ZN(n_648));
   NAND2_X1 i_698 (.A1(n_723), .A2(n_1743), .ZN(n_649));
   AOI22_X1 i_699 (.A1(b_mantissa[7]), .A2(a_mantissa[20]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[21]), .ZN(n_660));
   XOR2_X1 i_700 (.A(n_664), .B(n_663), .Z(n_1857));
   NAND2_X1 i_701 (.A1(b_mantissa[5]), .A2(a_mantissa[22]), .ZN(n_663));
   NAND2_X1 i_702 (.A1(n_667), .A2(n_665), .ZN(n_664));
   INV_X1 i_703 (.A(n_666), .ZN(n_665));
   AOI21_X1 i_704 (.A(b_mantissa[4]), .B1(b_mantissa[3]), .B2(n_724), .ZN(n_666));
   OAI211_X1 i_705 (.A(b_mantissa[4]), .B(n_736), .C1(n_1583), .C2(n_724), 
      .ZN(n_667));
   AOI21_X1 i_706 (.A(n_674), .B1(n_672), .B2(n_670), .ZN(n_1737));
   OAI21_X1 i_707 (.A(n_680), .B1(n_678), .B2(n_676), .ZN(n_1746));
   OAI21_X1 i_708 (.A(n_696), .B1(n_686), .B2(n_684), .ZN(n_1753));
   OAI21_X1 i_709 (.A(n_702), .B1(n_704), .B2(n_700), .ZN(n_1760));
   OAI21_X1 i_710 (.A(n_710), .B1(n_711), .B2(n_708), .ZN(n_1767));
   OAI21_X1 i_711 (.A(n_720), .B1(n_722), .B2(n_716), .ZN(n_1774));
   XOR2_X1 i_712 (.A(n_671), .B(n_670), .Z(n_1736));
   NAND2_X1 i_713 (.A1(b_mantissa[22]), .A2(a_mantissa[4]), .ZN(n_670));
   NAND2_X1 i_714 (.A1(n_673), .A2(n_672), .ZN(n_671));
   NAND3_X1 i_715 (.A1(b_mantissa[21]), .A2(a_mantissa[5]), .A3(a_mantissa[3]), 
      .ZN(n_672));
   INV_X1 i_716 (.A(n_674), .ZN(n_673));
   AOI21_X1 i_717 (.A(a_mantissa[3]), .B1(b_mantissa[21]), .B2(a_mantissa[5]), 
      .ZN(n_674));
   XNOR2_X1 i_718 (.A(n_677), .B(n_676), .ZN(n_1745));
   NAND2_X1 i_719 (.A1(b_mantissa[20]), .A2(a_mantissa[6]), .ZN(n_676));
   NOR2_X1 i_720 (.A1(n_679), .A2(n_678), .ZN(n_677));
   AOI21_X1 i_721 (.A(n_1635), .B1(b_mantissa[19]), .B2(a_mantissa[7]), .ZN(
      n_678));
   INV_X1 i_722 (.A(n_680), .ZN(n_679));
   NAND3_X1 i_723 (.A1(b_mantissa[19]), .A2(a_mantissa[7]), .A3(n_1635), 
      .ZN(n_680));
   XNOR2_X1 i_724 (.A(n_685), .B(n_684), .ZN(n_1752));
   NAND2_X1 i_725 (.A1(b_mantissa[17]), .A2(a_mantissa[9]), .ZN(n_684));
   NOR2_X1 i_726 (.A1(n_687), .A2(n_686), .ZN(n_685));
   AOI21_X1 i_727 (.A(n_1663), .B1(b_mantissa[16]), .B2(a_mantissa[10]), 
      .ZN(n_686));
   INV_X1 i_728 (.A(n_696), .ZN(n_687));
   NAND3_X1 i_729 (.A1(b_mantissa[16]), .A2(a_mantissa[10]), .A3(n_1663), 
      .ZN(n_696));
   XOR2_X1 i_730 (.A(n_701), .B(n_700), .Z(n_1759));
   NAND2_X1 i_731 (.A1(b_mantissa[14]), .A2(a_mantissa[12]), .ZN(n_700));
   NAND2_X1 i_732 (.A1(n_703), .A2(n_702), .ZN(n_701));
   NAND3_X1 i_733 (.A1(b_mantissa[13]), .A2(a_mantissa[13]), .A3(n_707), 
      .ZN(n_702));
   INV_X1 i_734 (.A(n_704), .ZN(n_703));
   AOI21_X1 i_735 (.A(n_707), .B1(b_mantissa[13]), .B2(a_mantissa[13]), .ZN(
      n_704));
   AND2_X1 i_736 (.A1(b_mantissa[12]), .A2(a_mantissa[14]), .ZN(n_707));
   XOR2_X1 i_737 (.A(n_709), .B(n_708), .Z(n_1766));
   NAND2_X1 i_738 (.A1(b_mantissa[11]), .A2(a_mantissa[15]), .ZN(n_708));
   NAND2_X1 i_739 (.A1(n_714), .A2(n_710), .ZN(n_709));
   OR3_X1 i_740 (.A1(n_554), .A2(n_957), .A3(n_715), .ZN(n_710));
   INV_X1 i_741 (.A(n_714), .ZN(n_711));
   OAI21_X1 i_742 (.A(n_715), .B1(n_554), .B2(n_957), .ZN(n_714));
   NAND2_X1 i_743 (.A1(b_mantissa[9]), .A2(a_mantissa[17]), .ZN(n_715));
   XOR2_X1 i_744 (.A(n_717), .B(n_716), .Z(n_1773));
   NAND2_X1 i_745 (.A1(b_mantissa[8]), .A2(a_mantissa[18]), .ZN(n_716));
   NAND2_X1 i_746 (.A1(n_721), .A2(n_720), .ZN(n_717));
   NAND3_X1 i_747 (.A1(b_mantissa[7]), .A2(a_mantissa[19]), .A3(n_723), .ZN(
      n_720));
   INV_X1 i_748 (.A(n_722), .ZN(n_721));
   AOI21_X1 i_749 (.A(n_723), .B1(b_mantissa[7]), .B2(a_mantissa[19]), .ZN(n_722));
   AND2_X1 i_750 (.A1(b_mantissa[6]), .A2(a_mantissa[20]), .ZN(n_723));
   XOR2_X1 i_751 (.A(n_735), .B(n_724), .Z(n_1779));
   AND2_X1 i_752 (.A1(b_mantissa[5]), .A2(a_mantissa[21]), .ZN(n_724));
   AOI21_X1 i_753 (.A(n_739), .B1(b_mantissa[4]), .B2(n_1583), .ZN(n_735));
   INV_X1 i_754 (.A(n_739), .ZN(n_736));
   AOI21_X1 i_755 (.A(b_mantissa[3]), .B1(b_mantissa[4]), .B2(a_mantissa[22]), 
      .ZN(n_739));
   OAI21_X1 i_756 (.A(n_750), .B1(n_753), .B2(n_748), .ZN(n_1668));
   OAI21_X1 i_757 (.A(n_756), .B1(n_759), .B2(n_754), .ZN(n_1675));
   OAI21_X1 i_758 (.A(n_762), .B1(n_776), .B2(n_760), .ZN(n_1682));
   OAI21_X1 i_759 (.A(n_781), .B1(n_783), .B2(n_779), .ZN(n_1689));
   OAI21_X1 i_760 (.A(n_788), .B1(n_790), .B2(n_786), .ZN(n_1696));
   NAND2_X1 i_761 (.A1(n_1584), .A2(n_740), .ZN(n_1703));
   NAND2_X1 i_762 (.A1(n_1585), .A2(n_1581), .ZN(n_740));
   XNOR2_X1 i_763 (.A(n_742), .B(n_1580), .ZN(n_1658));
   NOR2_X1 i_764 (.A1(n_1577), .A2(n_743), .ZN(n_742));
   INV_X1 i_765 (.A(n_1578), .ZN(n_743));
   XOR2_X1 i_766 (.A(n_749), .B(n_748), .Z(n_1667));
   NAND2_X1 i_767 (.A1(b_mantissa[20]), .A2(a_mantissa[5]), .ZN(n_748));
   NAND2_X1 i_768 (.A1(n_752), .A2(n_750), .ZN(n_749));
   NAND3_X1 i_769 (.A1(b_mantissa[18]), .A2(a_mantissa[7]), .A3(n_1430), 
      .ZN(n_750));
   INV_X1 i_770 (.A(n_753), .ZN(n_752));
   AOI21_X1 i_771 (.A(n_1430), .B1(b_mantissa[18]), .B2(a_mantissa[7]), .ZN(
      n_753));
   XOR2_X1 i_772 (.A(n_755), .B(n_754), .Z(n_1674));
   NAND2_X1 i_773 (.A1(b_mantissa[17]), .A2(a_mantissa[8]), .ZN(n_754));
   NAND2_X1 i_774 (.A1(n_757), .A2(n_756), .ZN(n_755));
   NAND3_X1 i_775 (.A1(b_mantissa[15]), .A2(a_mantissa[10]), .A3(n_1497), 
      .ZN(n_756));
   INV_X1 i_776 (.A(n_759), .ZN(n_757));
   AOI21_X1 i_777 (.A(n_1497), .B1(b_mantissa[15]), .B2(a_mantissa[10]), 
      .ZN(n_759));
   XOR2_X1 i_778 (.A(n_761), .B(n_760), .Z(n_1681));
   NAND2_X1 i_779 (.A1(b_mantissa[14]), .A2(a_mantissa[11]), .ZN(n_760));
   NAND2_X1 i_780 (.A1(n_775), .A2(n_762), .ZN(n_761));
   NAND3_X1 i_781 (.A1(b_mantissa[12]), .A2(a_mantissa[13]), .A3(n_1508), 
      .ZN(n_762));
   INV_X1 i_782 (.A(n_776), .ZN(n_775));
   AOI21_X1 i_783 (.A(n_1508), .B1(b_mantissa[12]), .B2(a_mantissa[13]), 
      .ZN(n_776));
   XOR2_X1 i_784 (.A(n_780), .B(n_779), .Z(n_1688));
   NAND2_X1 i_785 (.A1(b_mantissa[11]), .A2(a_mantissa[14]), .ZN(n_779));
   NAND2_X1 i_786 (.A1(n_782), .A2(n_781), .ZN(n_780));
   NAND3_X1 i_787 (.A1(b_mantissa[9]), .A2(a_mantissa[16]), .A3(n_1519), 
      .ZN(n_781));
   INV_X1 i_788 (.A(n_783), .ZN(n_782));
   AOI21_X1 i_789 (.A(n_1519), .B1(b_mantissa[9]), .B2(a_mantissa[16]), .ZN(
      n_783));
   XOR2_X1 i_790 (.A(n_787), .B(n_786), .Z(n_1695));
   NAND2_X1 i_791 (.A1(b_mantissa[8]), .A2(a_mantissa[17]), .ZN(n_786));
   NAND2_X1 i_792 (.A1(n_789), .A2(n_788), .ZN(n_787));
   NAND3_X1 i_793 (.A1(b_mantissa[6]), .A2(a_mantissa[19]), .A3(n_1449), 
      .ZN(n_788));
   INV_X1 i_794 (.A(n_790), .ZN(n_789));
   AOI21_X1 i_795 (.A(n_1449), .B1(b_mantissa[6]), .B2(a_mantissa[19]), .ZN(
      n_790));
   AOI21_X1 i_796 (.A(n_803), .B1(n_802), .B2(n_800), .ZN(n_1573));
   OAI21_X1 i_797 (.A(n_1429), .B1(n_1428), .B2(n_1427), .ZN(n_1582));
   XNOR2_X1 i_798 (.A(n_801), .B(n_800), .ZN(n_1572));
   NAND2_X1 i_799 (.A1(b_mantissa[22]), .A2(a_mantissa[2]), .ZN(n_800));
   AOI21_X1 i_800 (.A(n_803), .B1(a_mantissa[3]), .B2(n_1263), .ZN(n_801));
   NAND2_X1 i_801 (.A1(a_mantissa[3]), .A2(n_1263), .ZN(n_802));
   AOI21_X1 i_802 (.A(a_mantissa[1]), .B1(b_mantissa[21]), .B2(a_mantissa[3]), 
      .ZN(n_803));
   OAI22_X1 i_803 (.A1(n_1407), .A2(n_1223), .B1(n_893), .B2(n_891), .ZN(n_1487));
   OAI21_X1 i_804 (.A(n_897), .B1(n_899), .B2(n_894), .ZN(n_1496));
   OAI21_X1 i_805 (.A(n_902), .B1(n_905), .B2(n_900), .ZN(n_1503));
   OAI21_X1 i_806 (.A(n_924), .B1(n_928), .B2(n_906), .ZN(n_1510));
   XNOR2_X1 i_807 (.A(n_892), .B(n_891), .ZN(n_1486));
   NAND2_X1 i_808 (.A1(b_mantissa[22]), .A2(a_mantissa[1]), .ZN(n_891));
   AOI21_X1 i_809 (.A(n_893), .B1(a_mantissa[2]), .B2(n_1222), .ZN(n_892));
   AOI21_X1 i_810 (.A(a_mantissa[0]), .B1(b_mantissa[21]), .B2(a_mantissa[2]), 
      .ZN(n_893));
   XOR2_X1 i_811 (.A(n_895), .B(n_894), .Z(n_1495));
   NAND2_X1 i_812 (.A1(b_mantissa[20]), .A2(a_mantissa[3]), .ZN(n_894));
   NAND2_X1 i_813 (.A1(n_898), .A2(n_897), .ZN(n_895));
   NAND3_X1 i_814 (.A1(b_mantissa[19]), .A2(a_mantissa[4]), .A3(n_1333), 
      .ZN(n_897));
   INV_X1 i_815 (.A(n_899), .ZN(n_898));
   AOI21_X1 i_816 (.A(n_1333), .B1(b_mantissa[19]), .B2(a_mantissa[4]), .ZN(
      n_899));
   XOR2_X1 i_817 (.A(n_901), .B(n_900), .Z(n_1502));
   NAND2_X1 i_818 (.A1(b_mantissa[17]), .A2(a_mantissa[6]), .ZN(n_900));
   NAND2_X1 i_819 (.A1(n_904), .A2(n_902), .ZN(n_901));
   NAND3_X1 i_820 (.A1(b_mantissa[16]), .A2(a_mantissa[7]), .A3(n_1364), 
      .ZN(n_902));
   INV_X1 i_821 (.A(n_905), .ZN(n_904));
   AOI21_X1 i_822 (.A(n_1364), .B1(b_mantissa[16]), .B2(a_mantissa[7]), .ZN(
      n_905));
   XOR2_X1 i_823 (.A(n_907), .B(n_906), .Z(n_1509));
   NAND2_X1 i_824 (.A1(b_mantissa[14]), .A2(a_mantissa[9]), .ZN(n_906));
   NAND2_X1 i_825 (.A1(n_925), .A2(n_924), .ZN(n_907));
   NAND3_X1 i_826 (.A1(b_mantissa[13]), .A2(a_mantissa[10]), .A3(n_1380), 
      .ZN(n_924));
   INV_X1 i_827 (.A(n_928), .ZN(n_925));
   AOI21_X1 i_828 (.A(n_1380), .B1(b_mantissa[13]), .B2(a_mantissa[10]), 
      .ZN(n_928));
   XOR2_X1 i_829 (.A(n_930), .B(n_1594), .Z(n_1516));
   NAND2_X1 i_830 (.A1(n_932), .A2(n_1591), .ZN(n_930));
   INV_X1 i_831 (.A(n_1592), .ZN(n_932));
   XOR2_X1 i_832 (.A(n_937), .B(n_1601), .Z(n_1523));
   NAND2_X1 i_833 (.A1(n_939), .A2(n_1598), .ZN(n_937));
   INV_X1 i_834 (.A(n_1599), .ZN(n_939));
   XOR2_X1 i_835 (.A(n_944), .B(n_1608), .Z(n_1530));
   NAND2_X1 i_836 (.A1(n_946), .A2(n_1605), .ZN(n_944));
   INV_X1 i_837 (.A(n_1606), .ZN(n_946));
   XOR2_X1 i_838 (.A(n_951), .B(n_1489), .Z(n_1536));
   AOI21_X1 i_839 (.A(n_1476), .B1(b_mantissa[1]), .B2(n_1485), .ZN(n_951));
   AOI21_X1 i_840 (.A(n_1048), .B1(n_1049), .B2(n_1044), .ZN(n_1453));
   OAI21_X1 i_841 (.A(n_1260), .B1(n_1261), .B2(n_1259), .ZN(n_1405));
   OAI21_X1 i_842 (.A(n_1329), .B1(n_1326), .B2(n_1325), .ZN(n_1412));
   OAI21_X1 i_843 (.A(n_1360), .B1(n_1342), .B2(n_1334), .ZN(n_1419));
   OAI21_X1 i_844 (.A(n_1376), .B1(n_1374), .B2(n_1366), .ZN(n_1426));
   OAI21_X1 i_845 (.A(n_1268), .B1(n_1267), .B2(n_1266), .ZN(n_1433));
   OAI21_X1 i_846 (.A(n_1275), .B1(n_1274), .B2(n_1273), .ZN(n_1440));
   OAI21_X1 i_847 (.A(n_1292), .B1(n_1287), .B2(n_1280), .ZN(n_1447));
   XOR2_X1 i_848 (.A(n_1045), .B(n_1044), .Z(n_1452));
   NAND2_X1 i_849 (.A1(b_mantissa[1]), .A2(a_mantissa[21]), .ZN(n_1044));
   OAI21_X1 i_850 (.A(n_1049), .B1(n_1485), .B2(n_1050), .ZN(n_1045));
   NOR2_X1 i_851 (.A1(n_1485), .A2(n_1050), .ZN(n_1048));
   NAND2_X1 i_852 (.A1(n_1485), .A2(n_1050), .ZN(n_1049));
   AOI22_X1 i_853 (.A1(n_1147), .A2(n_1321), .B1(n_1134), .B2(n_1132), .ZN(
      n_1050));
   AOI21_X1 i_854 (.A(n_1058), .B1(n_1057), .B2(n_1055), .ZN(n_1373));
   OAI21_X1 i_855 (.A(n_1110), .B1(n_1112), .B2(n_1106), .ZN(n_1345));
   OAI21_X1 i_856 (.A(n_1118), .B1(n_1120), .B2(n_1114), .ZN(n_1352));
   OAI21_X1 i_857 (.A(n_1126), .B1(n_1128), .B2(n_1124), .ZN(n_1359));
   XNOR2_X1 i_858 (.A(n_1056), .B(n_1055), .ZN(n_1372));
   NAND2_X1 i_859 (.A1(b_mantissa[0]), .A2(a_mantissa[21]), .ZN(n_1055));
   AOI21_X1 i_860 (.A(n_1058), .B1(n_1062), .B2(n_1059), .ZN(n_1056));
   NAND2_X1 i_861 (.A1(n_1062), .A2(n_1059), .ZN(n_1057));
   NOR2_X1 i_862 (.A1(n_1062), .A2(n_1059), .ZN(n_1058));
   OAI21_X1 i_863 (.A(n_1195), .B1(n_1197), .B2(n_1191), .ZN(n_1059));
   OAI21_X1 i_864 (.A(n_1144), .B1(n_1156), .B2(n_1141), .ZN(n_1062));
   XOR2_X1 i_865 (.A(n_1065), .B(n_1223), .Z(n_1323));
   NAND2_X1 i_866 (.A1(n_1224), .A2(n_1066), .ZN(n_1065));
   INV_X1 i_867 (.A(n_1225), .ZN(n_1066));
   XOR2_X1 i_868 (.A(n_1073), .B(n_1229), .Z(n_1330));
   NAND2_X1 i_869 (.A1(n_1076), .A2(n_1233), .ZN(n_1073));
   INV_X1 i_870 (.A(n_1232), .ZN(n_1076));
   XOR2_X1 i_871 (.A(n_1080), .B(n_1234), .Z(n_1337));
   NAND2_X1 i_872 (.A1(n_1083), .A2(n_1248), .ZN(n_1080));
   INV_X1 i_873 (.A(n_1235), .ZN(n_1083));
   XOR2_X1 i_874 (.A(n_1107), .B(n_1106), .Z(n_1344));
   NAND2_X1 i_875 (.A1(b_mantissa[12]), .A2(a_mantissa[9]), .ZN(n_1106));
   NAND2_X1 i_876 (.A1(n_1111), .A2(n_1110), .ZN(n_1107));
   NAND3_X1 i_877 (.A1(b_mantissa[10]), .A2(a_mantissa[11]), .A3(n_1402), 
      .ZN(n_1110));
   INV_X1 i_878 (.A(n_1112), .ZN(n_1111));
   AOI21_X1 i_879 (.A(n_1402), .B1(b_mantissa[10]), .B2(a_mantissa[11]), 
      .ZN(n_1112));
   XOR2_X1 i_880 (.A(n_1117), .B(n_1114), .Z(n_1351));
   NAND2_X1 i_881 (.A1(b_mantissa[9]), .A2(a_mantissa[12]), .ZN(n_1114));
   NAND2_X1 i_882 (.A1(n_1119), .A2(n_1118), .ZN(n_1117));
   NAND3_X1 i_883 (.A1(b_mantissa[7]), .A2(a_mantissa[14]), .A3(n_1270), 
      .ZN(n_1118));
   INV_X1 i_884 (.A(n_1120), .ZN(n_1119));
   AOI21_X1 i_885 (.A(n_1270), .B1(b_mantissa[7]), .B2(a_mantissa[14]), .ZN(
      n_1120));
   XOR2_X1 i_886 (.A(n_1125), .B(n_1124), .Z(n_1358));
   NAND2_X1 i_887 (.A1(b_mantissa[6]), .A2(a_mantissa[15]), .ZN(n_1124));
   NAND2_X1 i_888 (.A1(n_1127), .A2(n_1126), .ZN(n_1125));
   NAND3_X1 i_889 (.A1(b_mantissa[4]), .A2(a_mantissa[17]), .A3(n_1277), 
      .ZN(n_1126));
   INV_X1 i_890 (.A(n_1128), .ZN(n_1127));
   AOI21_X1 i_891 (.A(n_1277), .B1(b_mantissa[4]), .B2(a_mantissa[17]), .ZN(
      n_1128));
   XNOR2_X1 i_892 (.A(n_1133), .B(n_1132), .ZN(n_1365));
   NAND2_X1 i_893 (.A1(b_mantissa[3]), .A2(a_mantissa[18]), .ZN(n_1132));
   AOI22_X1 i_894 (.A1(n_1145), .A2(n_1299), .B1(n_1147), .B2(n_1321), .ZN(
      n_1133));
   NAND2_X1 i_895 (.A1(n_1145), .A2(n_1299), .ZN(n_1134));
   OAI21_X1 i_896 (.A(n_1154), .B1(n_1176), .B2(n_1152), .ZN(n_1265));
   OAI21_X1 i_897 (.A(n_1181), .B1(n_1183), .B2(n_1177), .ZN(n_1272));
   OAI21_X1 i_898 (.A(n_1188), .B1(n_1190), .B2(n_1184), .ZN(n_1279));
   XOR2_X1 i_899 (.A(n_1140), .B(n_1249), .Z(n_1250));
   NAND2_X1 i_900 (.A1(n_1142), .A2(n_1253), .ZN(n_1140));
   INV_X1 i_901 (.A(n_1252), .ZN(n_1142));
   XOR2_X1 i_902 (.A(n_1146), .B(n_1254), .Z(n_1257));
   NAND2_X1 i_903 (.A1(n_1148), .A2(n_1256), .ZN(n_1146));
   INV_X1 i_904 (.A(n_1255), .ZN(n_1148));
   XOR2_X1 i_905 (.A(n_1153), .B(n_1152), .Z(n_1264));
   NAND2_X1 i_906 (.A1(b_mantissa[14]), .A2(a_mantissa[6]), .ZN(n_1152));
   NAND2_X1 i_907 (.A1(n_1155), .A2(n_1154), .ZN(n_1153));
   NAND3_X1 i_908 (.A1(b_mantissa[13]), .A2(a_mantissa[7]), .A3(n_1079), 
      .ZN(n_1154));
   INV_X1 i_909 (.A(n_1176), .ZN(n_1155));
   AOI21_X1 i_910 (.A(n_1079), .B1(b_mantissa[13]), .B2(a_mantissa[7]), .ZN(
      n_1176));
   XOR2_X1 i_911 (.A(n_1180), .B(n_1177), .Z(n_1271));
   NAND2_X1 i_912 (.A1(b_mantissa[11]), .A2(a_mantissa[9]), .ZN(n_1177));
   NAND2_X1 i_913 (.A1(n_1182), .A2(n_1181), .ZN(n_1180));
   NAND3_X1 i_914 (.A1(b_mantissa[10]), .A2(a_mantissa[10]), .A3(n_1087), 
      .ZN(n_1181));
   INV_X1 i_915 (.A(n_1183), .ZN(n_1182));
   AOI21_X1 i_916 (.A(n_1087), .B1(b_mantissa[10]), .B2(a_mantissa[10]), 
      .ZN(n_1183));
   XOR2_X1 i_917 (.A(n_1187), .B(n_1184), .Z(n_1278));
   NAND2_X1 i_918 (.A1(b_mantissa[8]), .A2(a_mantissa[12]), .ZN(n_1184));
   NAND2_X1 i_919 (.A1(n_1189), .A2(n_1188), .ZN(n_1187));
   NAND3_X1 i_920 (.A1(b_mantissa[7]), .A2(a_mantissa[13]), .A3(n_1131), 
      .ZN(n_1188));
   INV_X1 i_921 (.A(n_1190), .ZN(n_1189));
   AOI21_X1 i_922 (.A(n_1131), .B1(b_mantissa[7]), .B2(a_mantissa[13]), .ZN(
      n_1190));
   XOR2_X1 i_923 (.A(n_1194), .B(n_1191), .Z(n_1285));
   NAND2_X1 i_924 (.A1(b_mantissa[5]), .A2(a_mantissa[15]), .ZN(n_1191));
   NAND2_X1 i_925 (.A1(n_1196), .A2(n_1195), .ZN(n_1194));
   NAND3_X1 i_926 (.A1(b_mantissa[4]), .A2(a_mantissa[16]), .A3(n_1051), 
      .ZN(n_1195));
   INV_X1 i_927 (.A(n_1197), .ZN(n_1196));
   AOI21_X1 i_928 (.A(n_1051), .B1(b_mantissa[4]), .B2(a_mantissa[16]), .ZN(
      n_1197));
   AOI21_X1 i_929 (.A(n_1283), .B1(n_1284), .B2(n_1281), .ZN(n_1220));
   OAI21_X1 i_930 (.A(n_1085), .B1(n_1084), .B2(n_1082), .ZN(n_1200));
   OAI21_X1 i_931 (.A(n_1121), .B1(n_1113), .B2(n_1097), .ZN(n_1207));
   OAI21_X1 i_932 (.A(n_1037), .B1(n_1036), .B2(n_1033), .ZN(n_1214));
   XNOR2_X1 i_933 (.A(n_1282), .B(n_1281), .ZN(n_1219));
   NAND2_X1 i_934 (.A1(b_mantissa[1]), .A2(a_mantissa[18]), .ZN(n_1281));
   AOI21_X1 i_935 (.A(n_1283), .B1(n_1149), .B2(n_1286), .ZN(n_1282));
   NOR2_X1 i_936 (.A1(n_1149), .A2(n_1286), .ZN(n_1283));
   NAND2_X1 i_937 (.A1(n_1149), .A2(n_1286), .ZN(n_1284));
   AOI22_X1 i_938 (.A1(n_966), .A2(n_1063), .B1(n_1363), .B2(n_1361), .ZN(n_1286));
   AOI21_X1 i_939 (.A(n_1291), .B1(n_1290), .B2(n_1288), .ZN(n_1151));
   OAI21_X1 i_940 (.A(n_1339), .B1(n_1341), .B2(n_1335), .ZN(n_1123));
   OAI21_X1 i_941 (.A(n_1347), .B1(n_1349), .B2(n_1343), .ZN(n_1130));
   OAI21_X1 i_942 (.A(n_1355), .B1(n_1357), .B2(n_1353), .ZN(n_1137));
   XNOR2_X1 i_943 (.A(n_1289), .B(n_1288), .ZN(n_1150));
   NAND2_X1 i_944 (.A1(b_mantissa[0]), .A2(a_mantissa[18]), .ZN(n_1288));
   AOI21_X1 i_945 (.A(n_1291), .B1(n_1294), .B2(n_1293), .ZN(n_1289));
   NAND2_X1 i_946 (.A1(n_1294), .A2(n_1293), .ZN(n_1290));
   NOR2_X1 i_947 (.A1(n_1294), .A2(n_1293), .ZN(n_1291));
   OAI21_X1 i_948 (.A(n_1421), .B1(n_1423), .B2(n_1417), .ZN(n_1293));
   OAI21_X1 i_949 (.A(n_964), .B1(n_973), .B2(n_963), .ZN(n_1294));
   XOR2_X1 i_950 (.A(n_1296), .B(n_1004), .Z(n_1108));
   NAND2_X1 i_951 (.A1(n_1322), .A2(n_1008), .ZN(n_1296));
   INV_X1 i_952 (.A(n_1005), .ZN(n_1322));
   XOR2_X1 i_953 (.A(n_1328), .B(n_1009), .Z(n_1115));
   NAND2_X1 i_954 (.A1(n_1332), .A2(n_1011), .ZN(n_1328));
   INV_X1 i_955 (.A(n_1010), .ZN(n_1332));
   XOR2_X1 i_956 (.A(n_1336), .B(n_1335), .Z(n_1122));
   NAND2_X1 i_957 (.A1(b_mantissa[12]), .A2(a_mantissa[6]), .ZN(n_1335));
   NAND2_X1 i_958 (.A1(n_1340), .A2(n_1339), .ZN(n_1336));
   NAND3_X1 i_959 (.A1(b_mantissa[10]), .A2(a_mantissa[8]), .A3(n_1081), 
      .ZN(n_1339));
   INV_X1 i_960 (.A(n_1341), .ZN(n_1340));
   AOI21_X1 i_961 (.A(n_1081), .B1(b_mantissa[10]), .B2(a_mantissa[8]), .ZN(
      n_1341));
   XOR2_X1 i_962 (.A(n_1346), .B(n_1343), .Z(n_1129));
   NAND2_X1 i_963 (.A1(b_mantissa[9]), .A2(a_mantissa[9]), .ZN(n_1343));
   NAND2_X1 i_964 (.A1(n_1348), .A2(n_1347), .ZN(n_1346));
   NAND3_X1 i_965 (.A1(b_mantissa[7]), .A2(a_mantissa[11]), .A3(n_1096), 
      .ZN(n_1347));
   INV_X1 i_966 (.A(n_1349), .ZN(n_1348));
   AOI21_X1 i_967 (.A(n_1096), .B1(b_mantissa[7]), .B2(a_mantissa[11]), .ZN(
      n_1349));
   XOR2_X1 i_968 (.A(n_1354), .B(n_1353), .Z(n_1136));
   NAND2_X1 i_969 (.A1(b_mantissa[6]), .A2(a_mantissa[12]), .ZN(n_1353));
   NAND2_X1 i_970 (.A1(n_1356), .A2(n_1355), .ZN(n_1354));
   NAND3_X1 i_971 (.A1(b_mantissa[4]), .A2(a_mantissa[14]), .A3(n_1135), 
      .ZN(n_1355));
   INV_X1 i_972 (.A(n_1357), .ZN(n_1356));
   AOI21_X1 i_973 (.A(n_1135), .B1(b_mantissa[4]), .B2(a_mantissa[14]), .ZN(
      n_1357));
   XNOR2_X1 i_974 (.A(n_1362), .B(n_1361), .ZN(n_1143));
   NAND2_X1 i_975 (.A1(b_mantissa[3]), .A2(a_mantissa[15]), .ZN(n_1361));
   AOI22_X1 i_976 (.A1(n_965), .A2(n_1052), .B1(n_966), .B2(n_1063), .ZN(n_1362));
   NAND2_X1 i_977 (.A1(n_965), .A2(n_1052), .ZN(n_1363));
   OAI21_X1 i_978 (.A(n_1369), .B1(n_1371), .B2(n_1367), .ZN(n_1047));
   XOR2_X1 i_979 (.A(n_1368), .B(n_1367), .Z(n_1046));
   NAND2_X1 i_980 (.A1(b_mantissa[17]), .A2(a_mantissa[0]), .ZN(n_1367));
   NAND2_X1 i_981 (.A1(n_1370), .A2(n_1369), .ZN(n_1368));
   NAND3_X1 i_982 (.A1(b_mantissa[16]), .A2(a_mantissa[1]), .A3(n_795), .ZN(
      n_1369));
   INV_X1 i_983 (.A(n_1371), .ZN(n_1370));
   AOI21_X1 i_984 (.A(n_795), .B1(b_mantissa[16]), .B2(a_mantissa[1]), .ZN(
      n_1371));
   XOR2_X1 i_985 (.A(n_1375), .B(n_991), .Z(n_1053));
   NAND2_X1 i_986 (.A1(n_1377), .A2(n_995), .ZN(n_1375));
   INV_X1 i_987 (.A(n_994), .ZN(n_1377));
   XOR2_X1 i_988 (.A(n_1406), .B(n_996), .Z(n_1060));
   NAND2_X1 i_989 (.A1(n_1408), .A2(n_998), .ZN(n_1406));
   INV_X1 i_990 (.A(n_997), .ZN(n_1408));
   XOR2_X1 i_991 (.A(n_1413), .B(n_1001), .Z(n_1067));
   NAND2_X1 i_992 (.A1(n_1415), .A2(n_1003), .ZN(n_1413));
   INV_X1 i_993 (.A(n_1002), .ZN(n_1415));
   XOR2_X1 i_994 (.A(n_1420), .B(n_1417), .Z(n_1074));
   NAND2_X1 i_995 (.A1(b_mantissa[5]), .A2(a_mantissa[12]), .ZN(n_1417));
   NAND2_X1 i_996 (.A1(n_1422), .A2(n_1421), .ZN(n_1420));
   NAND3_X1 i_997 (.A1(b_mantissa[4]), .A2(a_mantissa[13]), .A3(n_953), .ZN(
      n_1421));
   INV_X1 i_998 (.A(n_1423), .ZN(n_1422));
   AOI21_X1 i_999 (.A(n_953), .B1(b_mantissa[4]), .B2(a_mantissa[13]), .ZN(
      n_1423));
   AOI21_X1 i_1000 (.A(n_936), .B1(n_1505), .B2(n_935), .ZN(n_1020));
   OAI21_X1 i_1001 (.A(n_794), .B1(n_796), .B2(n_763), .ZN(n_986));
   OAI21_X1 i_1002 (.A(n_804), .B1(n_799), .B2(n_797), .ZN(n_993));
   NAND2_X1 i_1003 (.A1(n_945), .A2(n_938), .ZN(n_1505));
   OAI21_X1 i_1004 (.A(n_1529), .B1(n_1533), .B2(n_1527), .ZN(n_934));
   OAI21_X1 i_1005 (.A(n_1538), .B1(n_1540), .B2(n_1535), .ZN(n_941));
   OAI21_X1 i_1006 (.A(n_1574), .B1(n_1576), .B2(n_1542), .ZN(n_948));
   XOR2_X1 i_1007 (.A(n_1520), .B(n_873), .Z(n_926));
   NAND2_X1 i_1008 (.A1(n_1522), .A2(n_877), .ZN(n_1520));
   INV_X1 i_1009 (.A(n_874), .ZN(n_1522));
   XOR2_X1 i_1010 (.A(n_1528), .B(n_1527), .Z(n_933));
   NAND2_X1 i_1011 (.A1(b_mantissa[12]), .A2(a_mantissa[3]), .ZN(n_1527));
   NAND2_X1 i_1012 (.A1(n_1532), .A2(n_1529), .ZN(n_1528));
   NAND3_X1 i_1013 (.A1(b_mantissa[10]), .A2(a_mantissa[5]), .A3(n_808), 
      .ZN(n_1529));
   INV_X1 i_1014 (.A(n_1533), .ZN(n_1532));
   AOI21_X1 i_1015 (.A(n_808), .B1(b_mantissa[10]), .B2(a_mantissa[5]), .ZN(
      n_1533));
   XOR2_X1 i_1016 (.A(n_1537), .B(n_1535), .Z(n_940));
   NAND2_X1 i_1017 (.A1(b_mantissa[9]), .A2(a_mantissa[6]), .ZN(n_1535));
   NAND2_X1 i_1018 (.A1(n_1539), .A2(n_1538), .ZN(n_1537));
   NAND3_X1 i_1019 (.A1(b_mantissa[7]), .A2(a_mantissa[8]), .A3(n_823), .ZN(
      n_1538));
   INV_X1 i_1020 (.A(n_1540), .ZN(n_1539));
   AOI21_X1 i_1021 (.A(n_823), .B1(b_mantissa[7]), .B2(a_mantissa[8]), .ZN(
      n_1540));
   XOR2_X1 i_1022 (.A(n_1571), .B(n_1542), .Z(n_947));
   NAND2_X1 i_1023 (.A1(b_mantissa[6]), .A2(a_mantissa[9]), .ZN(n_1542));
   NAND2_X1 i_1024 (.A1(n_1575), .A2(n_1574), .ZN(n_1571));
   NAND3_X1 i_1025 (.A1(b_mantissa[4]), .A2(a_mantissa[11]), .A3(n_950), 
      .ZN(n_1574));
   INV_X1 i_1026 (.A(n_1576), .ZN(n_1575));
   AOI21_X1 i_1027 (.A(n_950), .B1(b_mantissa[4]), .B2(a_mantissa[11]), .ZN(
      n_1576));
   XNOR2_X1 i_1028 (.A(n_1579), .B(n_943), .ZN(n_954));
   AOI22_X1 i_1029 (.A1(n_609), .A2(n_955), .B1(n_610), .B2(n_956), .ZN(n_1579));
   XOR2_X1 i_1030 (.A(n_1586), .B(n_851), .Z(n_875));
   NAND2_X1 i_1031 (.A1(n_1590), .A2(n_855), .ZN(n_1586));
   INV_X1 i_1032 (.A(n_854), .ZN(n_1590));
   XOR2_X1 i_1033 (.A(n_1593), .B(n_856), .Z(n_882));
   NAND2_X1 i_1034 (.A1(n_1597), .A2(n_858), .ZN(n_1593));
   INV_X1 i_1035 (.A(n_857), .ZN(n_1597));
   XOR2_X1 i_1036 (.A(n_1600), .B(n_859), .Z(n_889));
   NAND2_X1 i_1037 (.A1(n_1604), .A2(n_864), .ZN(n_1600));
   INV_X1 i_1038 (.A(n_863), .ZN(n_1604));
   XOR2_X1 i_1039 (.A(n_1607), .B(n_848), .Z(n_896));
   NAND2_X1 i_1040 (.A1(n_1611), .A2(n_850), .ZN(n_1607));
   INV_X1 i_1041 (.A(n_849), .ZN(n_1611));
   OAI21_X1 i_1042 (.A(n_588), .B1(n_587), .B2(n_586), .ZN(n_833));
   OAI21_X1 i_1043 (.A(n_596), .B1(n_595), .B2(n_594), .ZN(n_840));
   OAI21_X1 i_1044 (.A(n_562), .B1(n_561), .B2(n_559), .ZN(n_847));
   XNOR2_X1 i_1045 (.A(n_1685), .B(n_824), .ZN(n_852));
   AOI21_X1 i_1046 (.A(n_827), .B1(n_613), .B2(n_829), .ZN(n_1685));
   AOI21_X1 i_1047 (.A(n_1697), .B1(n_1694), .B2(n_1692), .ZN(n_806));
   XNOR2_X1 i_1048 (.A(n_1693), .B(n_1692), .ZN(n_805));
   NAND2_X1 i_1049 (.A1(b_mantissa[0]), .A2(a_mantissa[12]), .ZN(n_1692));
   AOI21_X1 i_1050 (.A(n_1697), .B1(n_1699), .B2(n_1698), .ZN(n_1693));
   NAND2_X1 i_1051 (.A1(n_1699), .A2(n_1698), .ZN(n_1694));
   NOR2_X1 i_1052 (.A1(n_1699), .A2(n_1698), .ZN(n_1697));
   OAI21_X1 i_1053 (.A(n_1777), .B1(n_1780), .B2(n_1775), .ZN(n_1698));
   OAI21_X1 i_1054 (.A(n_1783), .B1(n_1815), .B2(n_1781), .ZN(n_1699));
   XOR2_X1 i_1055 (.A(n_1701), .B(n_836), .Z(n_777));
   NAND2_X1 i_1056 (.A1(n_1705), .A2(n_838), .ZN(n_1701));
   INV_X1 i_1057 (.A(n_837), .ZN(n_1705));
   XOR2_X1 i_1058 (.A(n_1739), .B(n_841), .Z(n_784));
   NAND2_X1 i_1059 (.A1(n_1741), .A2(n_843), .ZN(n_1739));
   INV_X1 i_1060 (.A(n_842), .ZN(n_1741));
   XOR2_X1 i_1061 (.A(n_1747), .B(n_844), .Z(n_791));
   NAND2_X1 i_1062 (.A1(n_1749), .A2(n_846), .ZN(n_1747));
   INV_X1 i_1063 (.A(n_845), .ZN(n_1749));
   XNOR2_X1 i_1064 (.A(n_1755), .B(n_831), .ZN(n_798));
   AOI22_X1 i_1065 (.A1(n_834), .A2(n_564), .B1(n_835), .B2(n_565), .ZN(n_1755));
   XOR2_X1 i_1066 (.A(n_1762), .B(n_331), .Z(n_737));
   NAND2_X1 i_1067 (.A1(n_346), .A2(n_545), .ZN(n_1762));
   XOR2_X1 i_1068 (.A(n_1769), .B(n_546), .Z(n_744));
   NAND2_X1 i_1069 (.A1(n_1771), .A2(n_551), .ZN(n_1769));
   INV_X1 i_1070 (.A(n_547), .ZN(n_1771));
   XOR2_X1 i_1071 (.A(n_1776), .B(n_1775), .Z(n_751));
   NAND2_X1 i_1072 (.A1(b_mantissa[5]), .A2(a_mantissa[6]), .ZN(n_1775));
   NAND2_X1 i_1073 (.A1(n_1778), .A2(n_1777), .ZN(n_1776));
   NAND3_X1 i_1074 (.A1(b_mantissa[4]), .A2(a_mantissa[7]), .A3(n_327), .ZN(
      n_1777));
   INV_X1 i_1075 (.A(n_1780), .ZN(n_1778));
   AOI21_X1 i_1076 (.A(n_327), .B1(b_mantissa[4]), .B2(a_mantissa[7]), .ZN(
      n_1780));
   XOR2_X1 i_1077 (.A(n_1782), .B(n_1781), .Z(n_758));
   NAND2_X1 i_1078 (.A1(b_mantissa[2]), .A2(a_mantissa[9]), .ZN(n_1781));
   NAND2_X1 i_1079 (.A1(n_1812), .A2(n_1783), .ZN(n_1782));
   NAND2_X1 i_1080 (.A1(n_1847), .A2(n_834), .ZN(n_1783));
   INV_X1 i_1081 (.A(n_1815), .ZN(n_1812));
   AOI22_X1 i_1082 (.A1(b_mantissa[0]), .A2(a_mantissa[11]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[10]), .ZN(n_1815));
   AOI21_X1 i_1083 (.A(n_1845), .B1(n_1842), .B2(n_1840), .ZN(n_719));
   XOR2_X1 i_1084 (.A(n_1817), .B(n_309), .Z(n_698));
   NAND2_X1 i_1085 (.A1(n_1820), .A2(n_311), .ZN(n_1817));
   INV_X1 i_1086 (.A(n_310), .ZN(n_1820));
   XOR2_X1 i_1087 (.A(n_1825), .B(n_312), .Z(n_705));
   NAND2_X1 i_1088 (.A1(n_320), .A2(n_1826), .ZN(n_1825));
   INV_X1 i_1089 (.A(n_318), .ZN(n_1826));
   XOR2_X1 i_1090 (.A(n_1833), .B(n_323), .Z(n_712));
   NAND2_X1 i_1091 (.A1(n_326), .A2(n_1834), .ZN(n_1833));
   INV_X1 i_1092 (.A(n_325), .ZN(n_1834));
   XNOR2_X1 i_1093 (.A(n_1841), .B(n_1840), .ZN(n_718));
   NAND2_X1 i_1094 (.A1(b_mantissa[1]), .A2(a_mantissa[9]), .ZN(n_1840));
   AOI21_X1 i_1095 (.A(n_1845), .B1(n_1847), .B2(n_1846), .ZN(n_1841));
   NAND2_X1 i_1096 (.A1(n_1847), .A2(n_1846), .ZN(n_1842));
   NOR2_X1 i_1097 (.A1(n_1847), .A2(n_1846), .ZN(n_1845));
   AOI22_X1 i_1098 (.A1(n_1923), .A2(n_330), .B1(n_1899), .B2(n_1895), .ZN(
      n_1846));
   NOR2_X1 i_1099 (.A1(n_958), .A2(n_2100), .ZN(n_1847));
   AOI21_X1 i_1100 (.A(n_1853), .B1(n_1852), .B2(n_1848), .ZN(n_683));
   OAI21_X1 i_1101 (.A(n_1860), .B1(n_1862), .B2(n_1856), .ZN(n_662));
   OAI21_X1 i_1102 (.A(n_1891), .B1(n_1893), .B2(n_1887), .ZN(n_669));
   XNOR2_X1 i_1103 (.A(n_1849), .B(n_1848), .ZN(n_682));
   NAND2_X1 i_1104 (.A1(b_mantissa[0]), .A2(a_mantissa[9]), .ZN(n_1848));
   AOI21_X1 i_1105 (.A(n_1853), .B1(n_1855), .B2(n_1854), .ZN(n_1849));
   NAND2_X1 i_1106 (.A1(n_1855), .A2(n_1854), .ZN(n_1852));
   NOR2_X1 i_1107 (.A1(n_1855), .A2(n_1854), .ZN(n_1853));
   OAI21_X1 i_1108 (.A(n_1914), .B1(n_1916), .B2(n_1910), .ZN(n_1854));
   OAI21_X1 i_1109 (.A(n_1921), .B1(n_1927), .B2(n_1917), .ZN(n_1855));
   XOR2_X1 i_1110 (.A(n_1859), .B(n_1856), .Z(n_661));
   NAND2_X1 i_1111 (.A1(b_mantissa[9]), .A2(a_mantissa[0]), .ZN(n_1856));
   NAND2_X1 i_1112 (.A1(n_1861), .A2(n_1860), .ZN(n_1859));
   NAND3_X1 i_1113 (.A1(b_mantissa[8]), .A2(a_mantissa[1]), .A3(n_1907), 
      .ZN(n_1860));
   INV_X1 i_1114 (.A(n_1862), .ZN(n_1861));
   AOI21_X1 i_1115 (.A(n_1907), .B1(b_mantissa[8]), .B2(a_mantissa[1]), .ZN(
      n_1862));
   XOR2_X1 i_1116 (.A(n_1890), .B(n_1887), .Z(n_668));
   NAND2_X1 i_1117 (.A1(b_mantissa[6]), .A2(a_mantissa[3]), .ZN(n_1887));
   NAND2_X1 i_1118 (.A1(n_1892), .A2(n_1891), .ZN(n_1890));
   NAND3_X1 i_1119 (.A1(b_mantissa[4]), .A2(a_mantissa[5]), .A3(n_321), .ZN(
      n_1891));
   INV_X1 i_1120 (.A(n_1893), .ZN(n_1892));
   AOI21_X1 i_1121 (.A(n_321), .B1(b_mantissa[4]), .B2(a_mantissa[5]), .ZN(
      n_1893));
   XNOR2_X1 i_1122 (.A(n_1896), .B(n_1895), .ZN(n_675));
   NAND2_X1 i_1123 (.A1(b_mantissa[3]), .A2(a_mantissa[6]), .ZN(n_1895));
   AOI22_X1 i_1124 (.A1(n_1922), .A2(n_329), .B1(n_1923), .B2(n_330), .ZN(n_1896));
   NAND2_X1 i_1125 (.A1(n_1922), .A2(n_329), .ZN(n_1899));
   OAI21_X1 i_1126 (.A(n_1906), .B1(n_1909), .B2(n_1902), .ZN(n_633));
   XOR2_X1 i_1127 (.A(n_1903), .B(n_1902), .Z(n_632));
   NAND2_X1 i_1128 (.A1(b_mantissa[8]), .A2(a_mantissa[0]), .ZN(n_1902));
   NAND2_X1 i_1129 (.A1(n_1908), .A2(n_1906), .ZN(n_1903));
   NAND3_X1 i_1130 (.A1(b_mantissa[6]), .A2(a_mantissa[1]), .A3(n_1907), 
      .ZN(n_1906));
   NOR2_X1 i_1131 (.A1(n_1445), .A2(n_1407), .ZN(n_1907));
   INV_X1 i_1132 (.A(n_1909), .ZN(n_1908));
   AOI22_X1 i_1133 (.A1(b_mantissa[6]), .A2(a_mantissa[2]), .B1(b_mantissa[7]), 
      .B2(a_mantissa[1]), .ZN(n_1909));
   XOR2_X1 i_1134 (.A(n_1913), .B(n_1910), .Z(n_639));
   NAND2_X1 i_1135 (.A1(b_mantissa[5]), .A2(a_mantissa[3]), .ZN(n_1910));
   NAND2_X1 i_1136 (.A1(n_1915), .A2(n_1914), .ZN(n_1913));
   NAND3_X1 i_1137 (.A1(b_mantissa[4]), .A2(a_mantissa[4]), .A3(n_1967), 
      .ZN(n_1914));
   INV_X1 i_1138 (.A(n_1916), .ZN(n_1915));
   AOI21_X1 i_1139 (.A(n_1967), .B1(b_mantissa[4]), .B2(a_mantissa[4]), .ZN(
      n_1916));
   XOR2_X1 i_1140 (.A(n_1920), .B(n_1917), .Z(n_646));
   NAND2_X1 i_1141 (.A1(b_mantissa[2]), .A2(a_mantissa[6]), .ZN(n_1917));
   NAND2_X1 i_1142 (.A1(n_1924), .A2(n_1921), .ZN(n_1920));
   NAND2_X1 i_1143 (.A1(n_1974), .A2(n_1922), .ZN(n_1921));
   INV_X1 i_1144 (.A(n_1923), .ZN(n_1922));
   NAND2_X1 i_1145 (.A1(b_mantissa[1]), .A2(a_mantissa[8]), .ZN(n_1923));
   INV_X1 i_1146 (.A(n_1927), .ZN(n_1924));
   AOI22_X1 i_1147 (.A1(b_mantissa[0]), .A2(a_mantissa[8]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[7]), .ZN(n_1927));
   NAND2_X1 i_1148 (.A1(n_1969), .A2(n_1928), .ZN(n_618));
   NAND2_X1 i_1149 (.A1(n_1975), .A2(n_1970), .ZN(n_1928));
   OAI21_X1 i_1150 (.A(n_1957), .B1(n_1959), .B2(n_1929), .ZN(n_605));
   OAI21_X1 i_1151 (.A(n_1966), .B1(n_1963), .B2(n_1960), .ZN(n_612));
   XOR2_X1 i_1152 (.A(n_1954), .B(n_1929), .Z(n_604));
   NAND2_X1 i_1153 (.A1(b_mantissa[7]), .A2(a_mantissa[0]), .ZN(n_1929));
   NAND2_X1 i_1154 (.A1(n_1958), .A2(n_1957), .ZN(n_1954));
   NAND3_X1 i_1155 (.A1(b_mantissa[6]), .A2(a_mantissa[2]), .A3(n_1992), 
      .ZN(n_1957));
   INV_X1 i_1156 (.A(n_1959), .ZN(n_1958));
   AOI22_X1 i_1157 (.A1(b_mantissa[5]), .A2(a_mantissa[2]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[1]), .ZN(n_1959));
   XOR2_X1 i_1158 (.A(n_1961), .B(n_1960), .Z(n_611));
   NAND2_X1 i_1159 (.A1(b_mantissa[4]), .A2(a_mantissa[3]), .ZN(n_1960));
   NAND2_X1 i_1160 (.A1(n_1966), .A2(n_1962), .ZN(n_1961));
   INV_X1 i_1161 (.A(n_1963), .ZN(n_1962));
   AOI22_X1 i_1162 (.A1(b_mantissa[2]), .A2(a_mantissa[5]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[4]), .ZN(n_1963));
   NAND3_X1 i_1163 (.A1(b_mantissa[2]), .A2(a_mantissa[4]), .A3(n_1967), 
      .ZN(n_1966));
   AND2_X1 i_1164 (.A1(b_mantissa[3]), .A2(a_mantissa[5]), .ZN(n_1967));
   XNOR2_X1 i_1165 (.A(n_1975), .B(n_1968), .ZN(n_617));
   NAND2_X1 i_1166 (.A1(n_1970), .A2(n_1969), .ZN(n_1968));
   NAND2_X1 i_1167 (.A1(n_1974), .A2(n_1973), .ZN(n_1969));
   OR2_X1 i_1168 (.A1(n_1974), .A2(n_1973), .ZN(n_1970));
   OAI21_X1 i_1169 (.A(n_1997), .B1(n_1996), .B2(n_1993), .ZN(n_1973));
   AND2_X1 i_1170 (.A1(b_mantissa[0]), .A2(a_mantissa[7]), .ZN(n_1974));
   NOR2_X1 i_1171 (.A1(n_1475), .A2(n_1431), .ZN(n_1975));
   AOI21_X1 i_1172 (.A(n_1981), .B1(n_1980), .B2(n_1976), .ZN(n_593));
   OAI21_X1 i_1173 (.A(n_1988), .B1(n_1990), .B2(n_1984), .ZN(n_579));
   XNOR2_X1 i_1174 (.A(n_1977), .B(n_1976), .ZN(n_592));
   NAND2_X1 i_1175 (.A1(b_mantissa[0]), .A2(a_mantissa[6]), .ZN(n_1976));
   AOI21_X1 i_1176 (.A(n_1981), .B1(n_1983), .B2(n_1982), .ZN(n_1977));
   NAND2_X1 i_1177 (.A1(n_1983), .A2(n_1982), .ZN(n_1980));
   NOR2_X1 i_1178 (.A1(n_1983), .A2(n_1982), .ZN(n_1981));
   OAI21_X1 i_1179 (.A(n_2029), .B1(n_2033), .B2(n_2027), .ZN(n_1982));
   OAI21_X1 i_1180 (.A(n_2024), .B1(n_2026), .B2(n_2020), .ZN(n_1983));
   XOR2_X1 i_1181 (.A(n_1987), .B(n_1984), .Z(n_578));
   NAND2_X1 i_1182 (.A1(b_mantissa[6]), .A2(a_mantissa[0]), .ZN(n_1984));
   NAND2_X1 i_1183 (.A1(n_1989), .A2(n_1988), .ZN(n_1987));
   NAND3_X1 i_1184 (.A1(b_mantissa[4]), .A2(a_mantissa[2]), .A3(n_1992), 
      .ZN(n_1988));
   INV_X1 i_1185 (.A(n_1990), .ZN(n_1989));
   AOI21_X1 i_1186 (.A(n_1992), .B1(b_mantissa[4]), .B2(a_mantissa[2]), .ZN(
      n_1990));
   AND2_X1 i_1187 (.A1(b_mantissa[5]), .A2(a_mantissa[1]), .ZN(n_1992));
   XOR2_X1 i_1188 (.A(n_1994), .B(n_1993), .Z(n_585));
   NAND2_X1 i_1189 (.A1(b_mantissa[3]), .A2(a_mantissa[3]), .ZN(n_1993));
   NAND2_X1 i_1190 (.A1(n_1997), .A2(n_1995), .ZN(n_1994));
   INV_X1 i_1191 (.A(n_1996), .ZN(n_1995));
   AOI22_X1 i_1192 (.A1(b_mantissa[2]), .A2(a_mantissa[4]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[5]), .ZN(n_1996));
   NAND3_X1 i_1193 (.A1(b_mantissa[2]), .A2(a_mantissa[5]), .A3(n_2046), 
      .ZN(n_1997));
   XOR2_X1 i_1194 (.A(n_2023), .B(n_2020), .Z(n_560));
   NAND2_X1 i_1195 (.A1(b_mantissa[5]), .A2(a_mantissa[0]), .ZN(n_2020));
   NAND2_X1 i_1196 (.A1(n_2025), .A2(n_2024), .ZN(n_2023));
   NAND3_X1 i_1197 (.A1(b_mantissa[4]), .A2(a_mantissa[1]), .A3(n_2040), 
      .ZN(n_2024));
   INV_X1 i_1198 (.A(n_2026), .ZN(n_2025));
   AOI21_X1 i_1199 (.A(n_2040), .B1(b_mantissa[4]), .B2(a_mantissa[1]), .ZN(
      n_2026));
   XOR2_X1 i_1200 (.A(n_2028), .B(n_2027), .Z(n_567));
   NAND2_X1 i_1201 (.A1(b_mantissa[2]), .A2(a_mantissa[3]), .ZN(n_2027));
   NAND2_X1 i_1202 (.A1(n_2032), .A2(n_2029), .ZN(n_2028));
   NAND3_X1 i_1203 (.A1(b_mantissa[0]), .A2(a_mantissa[5]), .A3(n_2046), 
      .ZN(n_2029));
   INV_X1 i_1204 (.A(n_2033), .ZN(n_2032));
   AOI21_X1 i_1205 (.A(n_2046), .B1(b_mantissa[0]), .B2(a_mantissa[5]), .ZN(
      n_2033));
   AOI21_X1 i_1206 (.A(n_2036), .B1(n_2039), .B2(n_2034), .ZN(n_544));
   NAND2_X1 i_1207 (.A1(b_mantissa[4]), .A2(a_mantissa[0]), .ZN(n_2034));
   INV_X1 i_1208 (.A(n_2036), .ZN(n_2035));
   AOI22_X1 i_1209 (.A1(b_mantissa[2]), .A2(a_mantissa[2]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[1]), .ZN(n_2036));
   NAND3_X1 i_1210 (.A1(b_mantissa[2]), .A2(a_mantissa[1]), .A3(n_2040), 
      .ZN(n_2039));
   AND2_X1 i_1211 (.A1(b_mantissa[3]), .A2(a_mantissa[2]), .ZN(n_2040));
   OAI21_X1 i_1212 (.A(n_2042), .B1(n_550), .B2(n_2041), .ZN(n_549));
   NAND2_X1 i_1213 (.A1(b_mantissa[1]), .A2(a_mantissa[3]), .ZN(n_2041));
   NAND2_X1 i_1214 (.A1(a_mantissa[4]), .A2(n_2043), .ZN(n_2042));
   OAI22_X1 i_1215 (.A1(n_2088), .A2(n_2048), .B1(n_958), .B2(n_550), .ZN(n_2043));
   AOI21_X1 i_1216 (.A(n_2048), .B1(n_2088), .B2(n_2047), .ZN(n_550));
   INV_X1 i_1217 (.A(n_2047), .ZN(n_2046));
   NAND2_X1 i_1218 (.A1(b_mantissa[1]), .A2(a_mantissa[4]), .ZN(n_2047));
   NAND2_X1 i_1219 (.A1(b_mantissa[0]), .A2(a_mantissa[3]), .ZN(n_2048));
   OAI21_X1 i_1220 (.A(n_2056), .B1(n_2054), .B2(n_2049), .ZN(n_534));
   NAND2_X1 i_1221 (.A1(b_mantissa[3]), .A2(a_mantissa[0]), .ZN(n_2049));
   AND2_X1 i_1222 (.A1(n_2060), .A2(n_2050), .ZN(o_mantissa[1]));
   OAI22_X1 i_1223 (.A1(n_1475), .A2(n_2096), .B1(n_958), .B2(n_553), .ZN(n_2050));
   OAI22_X1 i_1224 (.A1(n_2061), .A2(n_2057), .B1(n_2060), .B2(n_2053), .ZN(
      o_mantissa[2]));
   NAND2_X1 i_1225 (.A1(n_2056), .A2(n_2055), .ZN(n_2053));
   INV_X1 i_1226 (.A(n_2055), .ZN(n_2054));
   OAI21_X1 i_1227 (.A(n_2090), .B1(n_1475), .B2(n_1407), .ZN(n_2055));
   NAND3_X1 i_1228 (.A1(b_mantissa[2]), .A2(a_mantissa[2]), .A3(n_2091), 
      .ZN(n_2056));
   OAI21_X1 i_1229 (.A(n_2060), .B1(n_2084), .B2(n_2063), .ZN(n_2057));
   NAND2_X1 i_1230 (.A1(n_2091), .A2(o_mantissa[0]), .ZN(n_2060));
   NOR2_X1 i_1231 (.A1(n_958), .A2(n_2096), .ZN(o_mantissa[0]));
   INV_X1 i_1232 (.A(n_2062), .ZN(n_2061));
   NAND2_X1 i_1233 (.A1(n_2084), .A2(n_2063), .ZN(n_2062));
   NAND2_X1 i_1234 (.A1(b_mantissa[0]), .A2(a_mantissa[2]), .ZN(n_2063));
   OR2_X1 i_1235 (.A1(n_2089), .A2(n_2087), .ZN(n_2084));
   AOI21_X1 i_1236 (.A(n_2091), .B1(b_mantissa[2]), .B2(a_mantissa[0]), .ZN(
      n_2087));
   INV_X1 i_1237 (.A(n_2089), .ZN(n_2088));
   NOR3_X1 i_1238 (.A1(n_1475), .A2(n_2096), .A3(n_2090), .ZN(n_2089));
   NAND2_X1 i_1239 (.A1(b_mantissa[2]), .A2(a_mantissa[1]), .ZN(n_2090));
   NOR2_X1 i_1240 (.A1(n_1475), .A2(n_553), .ZN(n_2091));
   OAI21_X1 i_1241 (.A(o_mantissa[47]), .B1(n_2093), .B2(n_2092), .ZN(
      o_mantissa[46]));
   NAND2_X1 i_1242 (.A1(n_2093), .A2(n_2092), .ZN(o_mantissa[47]));
   INV_X1 i_1243 (.A(n_188), .ZN(n_2092));
   INV_X1 i_1244 (.A(n_145), .ZN(n_2093));
   INV_X1 i_1245 (.A(a_mantissa[0]), .ZN(n_2096));
   INV_X1 i_1246 (.A(a_mantissa[10]), .ZN(n_2100));
   INV_X1 i_1247 (.A(a_mantissa[17]), .ZN(n_2106));
   INV_X1 i_1248 (.A(a_mantissa[21]), .ZN(n_2111));
   INV_X1 i_1249 (.A(b_mantissa[16]), .ZN(n_266));
   FA_X1 i_1250 (.A(n_713), .B(n_706), .CI(n_699), .CO(n_764), .S(n_304));
   FA_X1 i_1251 (.A(n_745), .B(n_738), .CI(n_764), .CO(n_307), .S(n_306));
   OAI21_X1 i_1252 (.A(n_311), .B1(n_310), .B2(n_309), .ZN(n_699));
   AOI21_X1 i_1253 (.A(n_318), .B1(n_320), .B2(n_312), .ZN(n_706));
   AOI21_X1 i_1254 (.A(n_325), .B1(n_326), .B2(n_323), .ZN(n_713));
   OAI21_X1 i_1255 (.A(n_545), .B1(n_358), .B2(n_331), .ZN(n_738));
   OAI21_X1 i_1256 (.A(n_551), .B1(n_547), .B2(n_546), .ZN(n_745));
   NAND2_X1 i_1257 (.A1(b_mantissa[10]), .A2(a_mantissa[0]), .ZN(n_309));
   AOI22_X1 i_1258 (.A1(b_mantissa[8]), .A2(a_mantissa[2]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[1]), .ZN(n_310));
   NAND4_X1 i_1259 (.A1(b_mantissa[8]), .A2(a_mantissa[2]), .A3(b_mantissa[9]), 
      .A4(a_mantissa[1]), .ZN(n_311));
   NAND2_X1 i_1260 (.A1(b_mantissa[7]), .A2(a_mantissa[3]), .ZN(n_312));
   AOI22_X1 i_1261 (.A1(b_mantissa[5]), .A2(a_mantissa[5]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[4]), .ZN(n_318));
   NAND3_X1 i_1262 (.A1(b_mantissa[6]), .A2(a_mantissa[5]), .A3(n_321), .ZN(
      n_320));
   AND2_X1 i_1263 (.A1(b_mantissa[5]), .A2(a_mantissa[4]), .ZN(n_321));
   NAND2_X1 i_1264 (.A1(b_mantissa[4]), .A2(a_mantissa[6]), .ZN(n_323));
   AOI22_X1 i_1265 (.A1(b_mantissa[2]), .A2(a_mantissa[8]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[7]), .ZN(n_325));
   NAND2_X1 i_1266 (.A1(n_329), .A2(n_327), .ZN(n_326));
   AND2_X1 i_1267 (.A1(b_mantissa[3]), .A2(a_mantissa[8]), .ZN(n_327));
   INV_X1 i_1268 (.A(n_330), .ZN(n_329));
   NAND2_X1 i_1269 (.A1(b_mantissa[2]), .A2(a_mantissa[7]), .ZN(n_330));
   NAND2_X1 i_1270 (.A1(b_mantissa[11]), .A2(a_mantissa[0]), .ZN(n_331));
   INV_X1 i_1271 (.A(n_358), .ZN(n_346));
   AOI22_X1 i_1272 (.A1(b_mantissa[9]), .A2(a_mantissa[2]), .B1(b_mantissa[10]), 
      .B2(a_mantissa[1]), .ZN(n_358));
   NAND4_X1 i_1273 (.A1(b_mantissa[9]), .A2(a_mantissa[2]), .A3(b_mantissa[10]), 
      .A4(a_mantissa[1]), .ZN(n_545));
   NAND2_X1 i_1274 (.A1(b_mantissa[8]), .A2(a_mantissa[3]), .ZN(n_546));
   AOI22_X1 i_1275 (.A1(b_mantissa[6]), .A2(a_mantissa[5]), .B1(b_mantissa[7]), 
      .B2(a_mantissa[4]), .ZN(n_547));
   NAND4_X1 i_1276 (.A1(b_mantissa[6]), .A2(a_mantissa[5]), .A3(b_mantissa[7]), 
      .A4(a_mantissa[4]), .ZN(n_551));
   INV_X1 i_1277 (.A(a_mantissa[1]), .ZN(n_553));
   INV_X1 i_1278 (.A(b_mantissa[10]), .ZN(n_554));
   XNOR2_X1 i_1279 (.A(n_559), .B(n_558), .ZN(n_555));
   AOI21_X1 i_1280 (.A(n_561), .B1(n_564), .B2(n_563), .ZN(n_558));
   NAND2_X1 i_1281 (.A1(b_mantissa[4]), .A2(a_mantissa[9]), .ZN(n_559));
   AOI22_X1 i_1282 (.A1(b_mantissa[2]), .A2(a_mantissa[11]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[10]), .ZN(n_561));
   NAND2_X1 i_1283 (.A1(n_564), .A2(n_563), .ZN(n_562));
   AND2_X1 i_1284 (.A1(b_mantissa[3]), .A2(a_mantissa[11]), .ZN(n_563));
   INV_X1 i_1285 (.A(n_565), .ZN(n_564));
   NAND2_X1 i_1286 (.A1(b_mantissa[2]), .A2(a_mantissa[10]), .ZN(n_565));
   FA_X1 i_1287 (.A(n_839), .B(n_832), .CI(n_825), .CO(n_568), .S(n_566));
   XNOR2_X1 i_1288 (.A(n_576), .B(n_569), .ZN(n_825));
   AOI21_X1 i_1289 (.A(n_583), .B1(n_581), .B2(n_580), .ZN(n_569));
   XNOR2_X1 i_1290 (.A(n_586), .B(n_570), .ZN(n_832));
   AOI21_X1 i_1291 (.A(n_587), .B1(n_591), .B2(n_590), .ZN(n_570));
   XNOR2_X1 i_1292 (.A(n_594), .B(n_571), .ZN(n_839));
   AOI21_X1 i_1293 (.A(n_595), .B1(n_602), .B2(n_597), .ZN(n_571));
   NAND2_X1 i_1294 (.A1(b_mantissa[13]), .A2(a_mantissa[0]), .ZN(n_576));
   NAND2_X1 i_1295 (.A1(n_581), .A2(n_580), .ZN(n_577));
   AND2_X1 i_1296 (.A1(b_mantissa[12]), .A2(a_mantissa[2]), .ZN(n_580));
   AND2_X1 i_1297 (.A1(b_mantissa[11]), .A2(a_mantissa[1]), .ZN(n_581));
   AOI22_X1 i_1298 (.A1(b_mantissa[11]), .A2(a_mantissa[2]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[1]), .ZN(n_583));
   NAND2_X1 i_1299 (.A1(b_mantissa[10]), .A2(a_mantissa[3]), .ZN(n_586));
   AOI22_X1 i_1300 (.A1(b_mantissa[8]), .A2(a_mantissa[5]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[4]), .ZN(n_587));
   NAND2_X1 i_1301 (.A1(n_591), .A2(n_590), .ZN(n_588));
   AND2_X1 i_1302 (.A1(b_mantissa[9]), .A2(a_mantissa[5]), .ZN(n_590));
   AND2_X1 i_1303 (.A1(b_mantissa[8]), .A2(a_mantissa[4]), .ZN(n_591));
   NAND2_X1 i_1304 (.A1(b_mantissa[7]), .A2(a_mantissa[6]), .ZN(n_594));
   AOI22_X1 i_1305 (.A1(b_mantissa[5]), .A2(a_mantissa[8]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[7]), .ZN(n_595));
   NAND2_X1 i_1306 (.A1(n_602), .A2(n_597), .ZN(n_596));
   AND2_X1 i_1307 (.A1(b_mantissa[6]), .A2(a_mantissa[8]), .ZN(n_597));
   AND2_X1 i_1308 (.A1(b_mantissa[5]), .A2(a_mantissa[7]), .ZN(n_602));
   XNOR2_X1 i_1309 (.A(n_607), .B(n_606), .ZN(n_603));
   AOI21_X1 i_1310 (.A(n_614), .B1(n_613), .B2(n_609), .ZN(n_606));
   NAND2_X1 i_1311 (.A1(b_mantissa[2]), .A2(a_mantissa[12]), .ZN(n_607));
   NAND2_X1 i_1312 (.A1(n_613), .A2(n_609), .ZN(n_608));
   INV_X1 i_1313 (.A(n_610), .ZN(n_609));
   NAND2_X1 i_1314 (.A1(b_mantissa[1]), .A2(a_mantissa[14]), .ZN(n_610));
   AND2_X1 i_1315 (.A1(b_mantissa[0]), .A2(a_mantissa[13]), .ZN(n_613));
   AOI22_X1 i_1316 (.A1(b_mantissa[0]), .A2(a_mantissa[14]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[13]), .ZN(n_614));
   FA_X1 i_1317 (.A(n_890), .B(n_883), .CI(n_876), .CO(n_968), .S(n_967));
   FA_X1 i_1318 (.A(n_927), .B(n_968), .CI(n_962), .CO(n_615), .S(n_1028));
   FA_X1 i_1319 (.A(n_792), .B(n_785), .CI(n_778), .CO(n_860), .S(n_616));
   FA_X1 i_1320 (.A(n_826), .B(n_860), .CI(n_853), .CO(n_911), .S(n_619));
   FA_X1 i_1321 (.A(n_911), .B(n_967), .CI(n_961), .CO(n_974), .S(n_620));
   FA_X1 i_1322 (.A(n_999), .B(n_992), .CI(n_985), .CO(n_621), .S(n_1032));
   FA_X1 i_1323 (.A(n_1028), .B(n_974), .CI(n_1032), .CO(n_623), .S(n_622));
   XNOR2_X1 i_1324 (.A(n_763), .B(n_635), .ZN(n_985));
   NOR2_X1 i_1325 (.A1(n_796), .A2(n_793), .ZN(n_635));
   XNOR2_X1 i_1326 (.A(n_797), .B(n_636), .ZN(n_992));
   AOI21_X1 i_1327 (.A(n_799), .B1(n_808), .B2(n_807), .ZN(n_636));
   XNOR2_X1 i_1328 (.A(n_809), .B(n_650), .ZN(n_999));
   AOI21_X1 i_1329 (.A(n_810), .B1(n_823), .B2(n_812), .ZN(n_650));
   XNOR2_X1 i_1330 (.A(n_681), .B(n_659), .ZN(n_961));
   AOI21_X1 i_1331 (.A(n_741), .B1(n_747), .B2(n_746), .ZN(n_659));
   OAI22_X1 i_1332 (.A1(n_878), .A2(n_828), .B1(n_827), .B2(n_824), .ZN(n_853));
   OAI21_X1 i_1333 (.A(n_838), .B1(n_837), .B2(n_836), .ZN(n_778));
   OAI21_X1 i_1334 (.A(n_843), .B1(n_842), .B2(n_841), .ZN(n_785));
   OAI21_X1 i_1335 (.A(n_846), .B1(n_845), .B2(n_844), .ZN(n_792));
   OAI21_X1 i_1336 (.A(n_577), .B1(n_583), .B2(n_576), .ZN(n_826));
   AOI21_X1 i_1337 (.A(n_741), .B1(n_697), .B2(n_681), .ZN(n_962));
   NAND2_X1 i_1338 (.A1(b_mantissa[0]), .A2(a_mantissa[15]), .ZN(n_681));
   NAND2_X1 i_1339 (.A1(n_747), .A2(n_746), .ZN(n_697));
   NOR2_X1 i_1340 (.A1(n_747), .A2(n_746), .ZN(n_741));
   OAI21_X1 i_1341 (.A(n_850), .B1(n_849), .B2(n_848), .ZN(n_746));
   OAI21_X1 i_1342 (.A(n_608), .B1(n_614), .B2(n_607), .ZN(n_747));
   OAI21_X1 i_1343 (.A(n_855), .B1(n_854), .B2(n_851), .ZN(n_876));
   OAI21_X1 i_1344 (.A(n_858), .B1(n_857), .B2(n_856), .ZN(n_883));
   OAI21_X1 i_1345 (.A(n_864), .B1(n_863), .B2(n_859), .ZN(n_890));
   AOI21_X1 i_1346 (.A(n_874), .B1(n_877), .B2(n_873), .ZN(n_927));
   NAND2_X1 i_1347 (.A1(b_mantissa[16]), .A2(a_mantissa[0]), .ZN(n_763));
   INV_X1 i_1348 (.A(n_794), .ZN(n_793));
   NAND3_X1 i_1349 (.A1(b_mantissa[14]), .A2(a_mantissa[1]), .A3(n_795), 
      .ZN(n_794));
   AND2_X1 i_1350 (.A1(b_mantissa[15]), .A2(a_mantissa[2]), .ZN(n_795));
   AOI22_X1 i_1351 (.A1(b_mantissa[14]), .A2(a_mantissa[2]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[1]), .ZN(n_796));
   NAND2_X1 i_1352 (.A1(b_mantissa[13]), .A2(a_mantissa[3]), .ZN(n_797));
   AOI22_X1 i_1353 (.A1(b_mantissa[11]), .A2(a_mantissa[5]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[4]), .ZN(n_799));
   NAND2_X1 i_1354 (.A1(n_808), .A2(n_807), .ZN(n_804));
   AND2_X1 i_1355 (.A1(b_mantissa[12]), .A2(a_mantissa[5]), .ZN(n_807));
   AND2_X1 i_1356 (.A1(b_mantissa[11]), .A2(a_mantissa[4]), .ZN(n_808));
   NAND2_X1 i_1357 (.A1(b_mantissa[10]), .A2(a_mantissa[6]), .ZN(n_809));
   AOI22_X1 i_1358 (.A1(b_mantissa[8]), .A2(a_mantissa[8]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[7]), .ZN(n_810));
   NAND2_X1 i_1359 (.A1(n_823), .A2(n_812), .ZN(n_811));
   AND2_X1 i_1360 (.A1(b_mantissa[9]), .A2(a_mantissa[8]), .ZN(n_812));
   AND2_X1 i_1361 (.A1(b_mantissa[8]), .A2(a_mantissa[7]), .ZN(n_823));
   NAND2_X1 i_1362 (.A1(b_mantissa[1]), .A2(a_mantissa[12]), .ZN(n_824));
   NOR2_X1 i_1363 (.A1(n_613), .A2(n_829), .ZN(n_827));
   INV_X1 i_1364 (.A(n_829), .ZN(n_828));
   AOI22_X1 i_1365 (.A1(n_831), .A2(n_830), .B1(n_565), .B2(n_835), .ZN(n_829));
   NAND2_X1 i_1366 (.A1(n_564), .A2(n_834), .ZN(n_830));
   NAND2_X1 i_1367 (.A1(b_mantissa[3]), .A2(a_mantissa[9]), .ZN(n_831));
   INV_X1 i_1368 (.A(n_835), .ZN(n_834));
   NAND2_X1 i_1369 (.A1(b_mantissa[1]), .A2(a_mantissa[11]), .ZN(n_835));
   NAND2_X1 i_1370 (.A1(b_mantissa[12]), .A2(a_mantissa[0]), .ZN(n_836));
   AOI21_X1 i_1371 (.A(n_581), .B1(b_mantissa[10]), .B2(a_mantissa[2]), .ZN(
      n_837));
   NAND3_X1 i_1372 (.A1(b_mantissa[10]), .A2(a_mantissa[2]), .A3(n_581), 
      .ZN(n_838));
   NAND2_X1 i_1373 (.A1(b_mantissa[9]), .A2(a_mantissa[3]), .ZN(n_841));
   AOI21_X1 i_1374 (.A(n_591), .B1(b_mantissa[7]), .B2(a_mantissa[5]), .ZN(n_842));
   NAND3_X1 i_1375 (.A1(b_mantissa[7]), .A2(a_mantissa[5]), .A3(n_591), .ZN(
      n_843));
   NAND2_X1 i_1376 (.A1(b_mantissa[6]), .A2(a_mantissa[6]), .ZN(n_844));
   AOI21_X1 i_1377 (.A(n_602), .B1(b_mantissa[4]), .B2(a_mantissa[8]), .ZN(n_845));
   NAND3_X1 i_1378 (.A1(b_mantissa[4]), .A2(a_mantissa[8]), .A3(n_602), .ZN(
      n_846));
   NAND2_X1 i_1379 (.A1(b_mantissa[5]), .A2(a_mantissa[9]), .ZN(n_848));
   AOI21_X1 i_1380 (.A(n_563), .B1(b_mantissa[4]), .B2(a_mantissa[10]), .ZN(
      n_849));
   NAND3_X1 i_1381 (.A1(b_mantissa[4]), .A2(a_mantissa[10]), .A3(n_563), 
      .ZN(n_850));
   NAND2_X1 i_1382 (.A1(b_mantissa[14]), .A2(a_mantissa[0]), .ZN(n_851));
   AOI21_X1 i_1383 (.A(n_580), .B1(b_mantissa[13]), .B2(a_mantissa[1]), .ZN(
      n_854));
   NAND3_X1 i_1384 (.A1(b_mantissa[13]), .A2(a_mantissa[1]), .A3(n_580), 
      .ZN(n_855));
   NAND2_X1 i_1385 (.A1(b_mantissa[11]), .A2(a_mantissa[3]), .ZN(n_856));
   AOI21_X1 i_1386 (.A(n_590), .B1(b_mantissa[10]), .B2(a_mantissa[4]), .ZN(
      n_857));
   NAND3_X1 i_1387 (.A1(b_mantissa[10]), .A2(a_mantissa[4]), .A3(n_590), 
      .ZN(n_858));
   NAND2_X1 i_1388 (.A1(b_mantissa[8]), .A2(a_mantissa[6]), .ZN(n_859));
   AOI21_X1 i_1389 (.A(n_597), .B1(b_mantissa[7]), .B2(a_mantissa[7]), .ZN(n_863));
   NAND3_X1 i_1390 (.A1(b_mantissa[7]), .A2(a_mantissa[7]), .A3(n_597), .ZN(
      n_864));
   NAND2_X1 i_1391 (.A1(b_mantissa[15]), .A2(a_mantissa[0]), .ZN(n_873));
   AOI22_X1 i_1392 (.A1(b_mantissa[14]), .A2(a_mantissa[1]), .B1(b_mantissa[13]), 
      .B2(a_mantissa[2]), .ZN(n_874));
   NAND4_X1 i_1393 (.A1(b_mantissa[13]), .A2(a_mantissa[1]), .A3(b_mantissa[14]), 
      .A4(a_mantissa[2]), .ZN(n_877));
   INV_X1 i_1394 (.A(n_613), .ZN(n_878));
   FA_X1 i_1395 (.A(n_1014), .B(n_1007), .CI(n_1000), .CO(n_879), .S(n_1086));
   FA_X1 i_1396 (.A(n_1019), .B(n_1013), .CI(n_1006), .CO(n_1031), .S(n_880));
   FA_X1 i_1397 (.A(n_1086), .B(n_621), .CI(n_1031), .CO(n_884), .S(n_881));
   XNOR2_X1 i_1398 (.A(n_888), .B(n_885), .ZN(n_1006));
   AOI21_X1 i_1399 (.A(n_910), .B1(n_950), .B2(n_949), .ZN(n_885));
   XNOR2_X1 i_1400 (.A(n_929), .B(n_886), .ZN(n_1013));
   AOI21_X1 i_1401 (.A(n_931), .B1(n_955), .B2(n_953), .ZN(n_886));
   XNOR2_X1 i_1402 (.A(n_935), .B(n_887), .ZN(n_1019));
   AOI21_X1 i_1403 (.A(n_936), .B1(n_945), .B2(n_938), .ZN(n_887));
   OAI21_X1 i_1404 (.A(n_811), .B1(n_810), .B2(n_809), .ZN(n_1000));
   AOI21_X1 i_1405 (.A(n_910), .B1(n_903), .B2(n_888), .ZN(n_1007));
   NAND2_X1 i_1406 (.A1(b_mantissa[7]), .A2(a_mantissa[9]), .ZN(n_888));
   NAND2_X1 i_1407 (.A1(n_950), .A2(n_949), .ZN(n_903));
   AOI22_X1 i_1408 (.A1(b_mantissa[5]), .A2(a_mantissa[11]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[10]), .ZN(n_910));
   OAI22_X1 i_1409 (.A1(n_956), .A2(n_952), .B1(n_931), .B2(n_929), .ZN(n_1014));
   NAND2_X1 i_1410 (.A1(b_mantissa[4]), .A2(a_mantissa[12]), .ZN(n_929));
   AOI22_X1 i_1411 (.A1(b_mantissa[2]), .A2(a_mantissa[14]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[13]), .ZN(n_931));
   NAND2_X1 i_1412 (.A1(b_mantissa[1]), .A2(a_mantissa[15]), .ZN(n_935));
   NOR2_X1 i_1413 (.A1(n_945), .A2(n_938), .ZN(n_936));
   AOI22_X1 i_1414 (.A1(n_943), .A2(n_942), .B1(n_610), .B2(n_956), .ZN(n_938));
   NAND2_X1 i_1415 (.A1(n_609), .A2(n_955), .ZN(n_942));
   NAND2_X1 i_1416 (.A1(b_mantissa[3]), .A2(a_mantissa[12]), .ZN(n_943));
   NOR2_X1 i_1417 (.A1(n_958), .A2(n_957), .ZN(n_945));
   AND2_X1 i_1418 (.A1(b_mantissa[6]), .A2(a_mantissa[11]), .ZN(n_949));
   AND2_X1 i_1419 (.A1(b_mantissa[5]), .A2(a_mantissa[10]), .ZN(n_950));
   INV_X1 i_1420 (.A(n_953), .ZN(n_952));
   AND2_X1 i_1421 (.A1(b_mantissa[3]), .A2(a_mantissa[14]), .ZN(n_953));
   INV_X1 i_1422 (.A(n_956), .ZN(n_955));
   NAND2_X1 i_1423 (.A1(b_mantissa[2]), .A2(a_mantissa[13]), .ZN(n_956));
   INV_X1 i_1424 (.A(a_mantissa[16]), .ZN(n_957));
   INV_X1 i_1425 (.A(b_mantissa[0]), .ZN(n_958));
   XNOR2_X1 i_1426 (.A(n_963), .B(n_960), .ZN(n_959));
   AOI21_X1 i_1427 (.A(n_973), .B1(n_945), .B2(n_965), .ZN(n_960));
   NAND2_X1 i_1428 (.A1(b_mantissa[2]), .A2(a_mantissa[15]), .ZN(n_963));
   NAND2_X1 i_1429 (.A1(n_945), .A2(n_965), .ZN(n_964));
   INV_X1 i_1430 (.A(n_966), .ZN(n_965));
   NAND2_X1 i_1431 (.A1(b_mantissa[1]), .A2(a_mantissa[17]), .ZN(n_966));
   AOI22_X1 i_1432 (.A1(b_mantissa[0]), .A2(a_mantissa[17]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[16]), .ZN(n_973));
   FA_X1 i_1433 (.A(n_1068), .B(n_1061), .CI(n_1054), .CO(n_1157), .S(n_983));
   FA_X1 i_1434 (.A(n_1116), .B(n_1109), .CI(n_1157), .CO(n_984), .S(n_1228));
   FA_X1 i_1435 (.A(n_1185), .B(n_1178), .CI(n_1228), .CO(n_988), .S(n_987));
   OAI21_X1 i_1436 (.A(n_995), .B1(n_994), .B2(n_991), .ZN(n_1054));
   OAI21_X1 i_1437 (.A(n_998), .B1(n_997), .B2(n_996), .ZN(n_1061));
   OAI21_X1 i_1438 (.A(n_1003), .B1(n_1002), .B2(n_1001), .ZN(n_1068));
   OAI21_X1 i_1439 (.A(n_1008), .B1(n_1005), .B2(n_1004), .ZN(n_1109));
   AOI21_X1 i_1440 (.A(n_1010), .B1(n_1011), .B2(n_1009), .ZN(n_1116));
   XNOR2_X1 i_1441 (.A(n_1012), .B(n_989), .ZN(n_1178));
   NOR2_X1 i_1442 (.A1(n_1018), .A2(n_1015), .ZN(n_989));
   XNOR2_X1 i_1443 (.A(n_1021), .B(n_990), .ZN(n_1185));
   NOR2_X1 i_1444 (.A1(n_1023), .A2(n_1022), .ZN(n_990));
   NAND2_X1 i_1445 (.A1(b_mantissa[14]), .A2(a_mantissa[3]), .ZN(n_991));
   AOI21_X1 i_1446 (.A(n_807), .B1(b_mantissa[13]), .B2(a_mantissa[4]), .ZN(
      n_994));
   NAND3_X1 i_1447 (.A1(b_mantissa[13]), .A2(a_mantissa[4]), .A3(n_807), 
      .ZN(n_995));
   NAND2_X1 i_1448 (.A1(b_mantissa[11]), .A2(a_mantissa[6]), .ZN(n_996));
   AOI21_X1 i_1449 (.A(n_812), .B1(b_mantissa[10]), .B2(a_mantissa[7]), .ZN(
      n_997));
   NAND3_X1 i_1450 (.A1(b_mantissa[10]), .A2(a_mantissa[7]), .A3(n_812), 
      .ZN(n_998));
   NAND2_X1 i_1451 (.A1(b_mantissa[8]), .A2(a_mantissa[9]), .ZN(n_1001));
   AOI21_X1 i_1452 (.A(n_949), .B1(b_mantissa[7]), .B2(a_mantissa[10]), .ZN(
      n_1002));
   NAND3_X1 i_1453 (.A1(b_mantissa[7]), .A2(a_mantissa[10]), .A3(n_949), 
      .ZN(n_1003));
   NAND2_X1 i_1454 (.A1(b_mantissa[18]), .A2(a_mantissa[0]), .ZN(n_1004));
   AOI22_X1 i_1455 (.A1(b_mantissa[17]), .A2(a_mantissa[1]), .B1(b_mantissa[16]), 
      .B2(a_mantissa[2]), .ZN(n_1005));
   NAND4_X1 i_1456 (.A1(b_mantissa[17]), .A2(a_mantissa[1]), .A3(b_mantissa[16]), 
      .A4(a_mantissa[2]), .ZN(n_1008));
   NAND2_X1 i_1457 (.A1(b_mantissa[15]), .A2(a_mantissa[3]), .ZN(n_1009));
   AOI22_X1 i_1458 (.A1(b_mantissa[14]), .A2(a_mantissa[4]), .B1(b_mantissa[13]), 
      .B2(a_mantissa[5]), .ZN(n_1010));
   NAND4_X1 i_1459 (.A1(b_mantissa[14]), .A2(a_mantissa[5]), .A3(b_mantissa[13]), 
      .A4(a_mantissa[4]), .ZN(n_1011));
   NAND2_X1 i_1460 (.A1(b_mantissa[19]), .A2(a_mantissa[0]), .ZN(n_1012));
   INV_X1 i_1461 (.A(n_1016), .ZN(n_1015));
   NAND3_X1 i_1462 (.A1(b_mantissa[17]), .A2(a_mantissa[1]), .A3(n_1017), 
      .ZN(n_1016));
   AND2_X1 i_1463 (.A1(b_mantissa[18]), .A2(a_mantissa[2]), .ZN(n_1017));
   AOI22_X1 i_1464 (.A1(b_mantissa[17]), .A2(a_mantissa[2]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[1]), .ZN(n_1018));
   NAND2_X1 i_1465 (.A1(b_mantissa[16]), .A2(a_mantissa[3]), .ZN(n_1021));
   AOI22_X1 i_1466 (.A1(b_mantissa[14]), .A2(a_mantissa[5]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[4]), .ZN(n_1022));
   INV_X1 i_1467 (.A(n_1024), .ZN(n_1023));
   NAND3_X1 i_1468 (.A1(b_mantissa[14]), .A2(a_mantissa[4]), .A3(n_1025), 
      .ZN(n_1024));
   AND2_X1 i_1469 (.A1(b_mantissa[15]), .A2(a_mantissa[5]), .ZN(n_1025));
   XNOR2_X1 i_1470 (.A(n_1033), .B(n_1030), .ZN(n_1029));
   AOI21_X1 i_1471 (.A(n_1036), .B1(n_1052), .B2(n_1051), .ZN(n_1030));
   NAND2_X1 i_1472 (.A1(b_mantissa[4]), .A2(a_mantissa[15]), .ZN(n_1033));
   AOI22_X1 i_1473 (.A1(b_mantissa[2]), .A2(a_mantissa[17]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[16]), .ZN(n_1036));
   NAND2_X1 i_1474 (.A1(n_1052), .A2(n_1051), .ZN(n_1037));
   AND2_X1 i_1475 (.A1(b_mantissa[3]), .A2(a_mantissa[17]), .ZN(n_1051));
   INV_X1 i_1476 (.A(n_1063), .ZN(n_1052));
   NAND2_X1 i_1477 (.A1(b_mantissa[2]), .A2(a_mantissa[16]), .ZN(n_1063));
   FA_X1 i_1478 (.A(n_1206), .B(n_1199), .CI(n_1192), .CO(n_1069), .S(n_1064));
   XNOR2_X1 i_1479 (.A(n_1075), .B(n_1070), .ZN(n_1192));
   AOI21_X1 i_1480 (.A(n_1077), .B1(n_1081), .B2(n_1079), .ZN(n_1070));
   XNOR2_X1 i_1481 (.A(n_1082), .B(n_1071), .ZN(n_1199));
   AOI21_X1 i_1482 (.A(n_1084), .B1(n_1096), .B2(n_1087), .ZN(n_1071));
   XNOR2_X1 i_1483 (.A(n_1097), .B(n_1072), .ZN(n_1206));
   AOI21_X1 i_1484 (.A(n_1113), .B1(n_1135), .B2(n_1131), .ZN(n_1072));
   NAND2_X1 i_1485 (.A1(b_mantissa[13]), .A2(a_mantissa[6]), .ZN(n_1075));
   AOI22_X1 i_1486 (.A1(b_mantissa[11]), .A2(a_mantissa[8]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[7]), .ZN(n_1077));
   NAND2_X1 i_1487 (.A1(n_1081), .A2(n_1079), .ZN(n_1078));
   AND2_X1 i_1488 (.A1(b_mantissa[12]), .A2(a_mantissa[8]), .ZN(n_1079));
   AND2_X1 i_1489 (.A1(b_mantissa[11]), .A2(a_mantissa[7]), .ZN(n_1081));
   NAND2_X1 i_1490 (.A1(b_mantissa[10]), .A2(a_mantissa[9]), .ZN(n_1082));
   AOI22_X1 i_1491 (.A1(b_mantissa[8]), .A2(a_mantissa[11]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[10]), .ZN(n_1084));
   NAND2_X1 i_1492 (.A1(n_1096), .A2(n_1087), .ZN(n_1085));
   AND2_X1 i_1493 (.A1(b_mantissa[9]), .A2(a_mantissa[11]), .ZN(n_1087));
   AND2_X1 i_1494 (.A1(b_mantissa[8]), .A2(a_mantissa[10]), .ZN(n_1096));
   NAND2_X1 i_1495 (.A1(b_mantissa[7]), .A2(a_mantissa[12]), .ZN(n_1097));
   AOI22_X1 i_1496 (.A1(b_mantissa[5]), .A2(a_mantissa[14]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[13]), .ZN(n_1113));
   NAND2_X1 i_1497 (.A1(n_1135), .A2(n_1131), .ZN(n_1121));
   AND2_X1 i_1498 (.A1(b_mantissa[6]), .A2(a_mantissa[14]), .ZN(n_1131));
   AND2_X1 i_1499 (.A1(b_mantissa[5]), .A2(a_mantissa[13]), .ZN(n_1135));
   XNOR2_X1 i_1500 (.A(n_1141), .B(n_1139), .ZN(n_1138));
   AOI21_X1 i_1501 (.A(n_1156), .B1(n_1149), .B2(n_1145), .ZN(n_1139));
   NAND2_X1 i_1502 (.A1(b_mantissa[2]), .A2(a_mantissa[18]), .ZN(n_1141));
   NAND2_X1 i_1503 (.A1(n_1149), .A2(n_1145), .ZN(n_1144));
   INV_X1 i_1504 (.A(n_1147), .ZN(n_1145));
   NAND2_X1 i_1505 (.A1(b_mantissa[1]), .A2(a_mantissa[20]), .ZN(n_1147));
   NOR2_X1 i_1506 (.A1(n_1198), .A2(n_958), .ZN(n_1149));
   AOI22_X1 i_1507 (.A1(b_mantissa[0]), .A2(a_mantissa[20]), .B1(b_mantissa[1]), 
      .B2(a_mantissa[19]), .ZN(n_1156));
   INV_X1 i_1508 (.A(a_mantissa[19]), .ZN(n_1198));
   FA_X1 i_1509 (.A(n_1425), .B(n_1418), .CI(n_1411), .CO(n_1201), .S(n_1467));
   FA_X1 i_1510 (.A(n_1446), .B(n_1439), .CI(n_1432), .CO(n_1202), .S(n_1465));
   FA_X1 i_1511 (.A(n_1193), .B(n_1186), .CI(n_1179), .CO(n_1300), .S(n_1203));
   FA_X1 i_1512 (.A(n_1258), .B(n_1251), .CI(n_1300), .CO(n_1381), .S(n_1204));
   FA_X1 i_1513 (.A(n_1338), .B(n_1331), .CI(n_1324), .CO(n_1205), .S(n_1461));
   FA_X1 i_1514 (.A(n_1404), .B(n_1381), .CI(n_1461), .CO(n_1208), .S(n_1469));
   FA_X1 i_1515 (.A(n_1467), .B(n_1465), .CI(n_1469), .CO(n_1210), .S(n_1209));
   INV_X1 i_1516 (.A(n_1211), .ZN(n_1324));
   OAI21_X1 i_1517 (.A(n_1224), .B1(n_1225), .B2(n_1222), .ZN(n_1211));
   AOI21_X1 i_1518 (.A(n_1232), .B1(n_1233), .B2(n_1229), .ZN(n_1331));
   OAI21_X1 i_1519 (.A(n_1248), .B1(n_1235), .B2(n_1234), .ZN(n_1338));
   OAI21_X1 i_1520 (.A(n_1016), .B1(n_1018), .B2(n_1012), .ZN(n_1179));
   OAI21_X1 i_1521 (.A(n_1024), .B1(n_1022), .B2(n_1021), .ZN(n_1186));
   OAI21_X1 i_1522 (.A(n_1078), .B1(n_1077), .B2(n_1075), .ZN(n_1193));
   OAI21_X1 i_1523 (.A(n_1253), .B1(n_1252), .B2(n_1249), .ZN(n_1251));
   OAI21_X1 i_1524 (.A(n_1256), .B1(n_1255), .B2(n_1254), .ZN(n_1258));
   XNOR2_X1 i_1525 (.A(n_1259), .B(n_1212), .ZN(n_1404));
   AOI21_X1 i_1526 (.A(n_1261), .B1(n_1263), .B2(n_1262), .ZN(n_1212));
   XNOR2_X1 i_1527 (.A(n_1266), .B(n_1213), .ZN(n_1432));
   AOI21_X1 i_1528 (.A(n_1267), .B1(n_1270), .B2(n_1269), .ZN(n_1213));
   XNOR2_X1 i_1529 (.A(n_1273), .B(n_1215), .ZN(n_1439));
   AOI21_X1 i_1530 (.A(n_1274), .B1(n_1277), .B2(n_1276), .ZN(n_1215));
   XNOR2_X1 i_1531 (.A(n_1280), .B(n_1216), .ZN(n_1446));
   AOI21_X1 i_1532 (.A(n_1287), .B1(n_1299), .B2(n_1295), .ZN(n_1216));
   XNOR2_X1 i_1533 (.A(n_1325), .B(n_1217), .ZN(n_1411));
   NOR2_X1 i_1534 (.A1(n_1327), .A2(n_1326), .ZN(n_1217));
   XNOR2_X1 i_1535 (.A(n_1334), .B(n_1218), .ZN(n_1418));
   NOR2_X1 i_1536 (.A1(n_1350), .A2(n_1342), .ZN(n_1218));
   XNOR2_X1 i_1537 (.A(n_1366), .B(n_1221), .ZN(n_1425));
   AOI21_X1 i_1538 (.A(n_1374), .B1(n_1402), .B2(n_1380), .ZN(n_1221));
   INV_X1 i_1539 (.A(n_1223), .ZN(n_1222));
   NAND2_X1 i_1540 (.A1(b_mantissa[21]), .A2(a_mantissa[0]), .ZN(n_1223));
   OAI22_X1 i_1541 (.A1(n_1410), .A2(n_1403), .B1(n_1409), .B2(n_1407), .ZN(
      n_1224));
   AND3_X1 i_1542 (.A1(b_mantissa[19]), .A2(a_mantissa[1]), .A3(n_1262), 
      .ZN(n_1225));
   NAND2_X1 i_1543 (.A1(b_mantissa[18]), .A2(a_mantissa[3]), .ZN(n_1229));
   AOI22_X1 i_1544 (.A1(b_mantissa[17]), .A2(a_mantissa[4]), .B1(b_mantissa[16]), 
      .B2(a_mantissa[5]), .ZN(n_1232));
   NAND4_X1 i_1545 (.A1(b_mantissa[17]), .A2(a_mantissa[5]), .A3(b_mantissa[16]), 
      .A4(a_mantissa[4]), .ZN(n_1233));
   NAND2_X1 i_1546 (.A1(b_mantissa[15]), .A2(a_mantissa[6]), .ZN(n_1234));
   AOI22_X1 i_1547 (.A1(b_mantissa[14]), .A2(a_mantissa[7]), .B1(b_mantissa[13]), 
      .B2(a_mantissa[8]), .ZN(n_1235));
   NAND4_X1 i_1548 (.A1(b_mantissa[14]), .A2(a_mantissa[7]), .A3(b_mantissa[13]), 
      .A4(a_mantissa[8]), .ZN(n_1248));
   NAND2_X1 i_1549 (.A1(b_mantissa[20]), .A2(a_mantissa[0]), .ZN(n_1249));
   AOI21_X1 i_1550 (.A(n_1017), .B1(b_mantissa[19]), .B2(a_mantissa[1]), 
      .ZN(n_1252));
   NAND3_X1 i_1551 (.A1(b_mantissa[19]), .A2(a_mantissa[1]), .A3(n_1017), 
      .ZN(n_1253));
   NAND2_X1 i_1552 (.A1(b_mantissa[17]), .A2(a_mantissa[3]), .ZN(n_1254));
   AOI21_X1 i_1553 (.A(n_1025), .B1(b_mantissa[16]), .B2(a_mantissa[4]), 
      .ZN(n_1255));
   NAND3_X1 i_1554 (.A1(b_mantissa[16]), .A2(a_mantissa[4]), .A3(n_1025), 
      .ZN(n_1256));
   NAND2_X1 i_1555 (.A1(b_mantissa[22]), .A2(a_mantissa[0]), .ZN(n_1259));
   NAND2_X1 i_1556 (.A1(n_1263), .A2(n_1262), .ZN(n_1260));
   NOR2_X1 i_1557 (.A1(n_1263), .A2(n_1262), .ZN(n_1261));
   NOR2_X1 i_1558 (.A1(n_1410), .A2(n_1407), .ZN(n_1262));
   NOR2_X1 i_1559 (.A1(n_1414), .A2(n_553), .ZN(n_1263));
   NAND2_X1 i_1560 (.A1(b_mantissa[10]), .A2(a_mantissa[12]), .ZN(n_1266));
   AOI22_X1 i_1561 (.A1(b_mantissa[8]), .A2(a_mantissa[14]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[13]), .ZN(n_1267));
   NAND2_X1 i_1562 (.A1(n_1270), .A2(n_1269), .ZN(n_1268));
   AND2_X1 i_1563 (.A1(b_mantissa[9]), .A2(a_mantissa[14]), .ZN(n_1269));
   AND2_X1 i_1564 (.A1(b_mantissa[8]), .A2(a_mantissa[13]), .ZN(n_1270));
   NAND2_X1 i_1565 (.A1(b_mantissa[7]), .A2(a_mantissa[15]), .ZN(n_1273));
   AOI22_X1 i_1566 (.A1(b_mantissa[5]), .A2(a_mantissa[17]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[16]), .ZN(n_1274));
   NAND2_X1 i_1567 (.A1(n_1277), .A2(n_1276), .ZN(n_1275));
   AND2_X1 i_1568 (.A1(b_mantissa[6]), .A2(a_mantissa[17]), .ZN(n_1276));
   AND2_X1 i_1569 (.A1(b_mantissa[5]), .A2(a_mantissa[16]), .ZN(n_1277));
   NAND2_X1 i_1570 (.A1(b_mantissa[4]), .A2(a_mantissa[18]), .ZN(n_1280));
   AOI22_X1 i_1571 (.A1(b_mantissa[2]), .A2(a_mantissa[20]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[19]), .ZN(n_1287));
   NAND2_X1 i_1572 (.A1(n_1299), .A2(n_1295), .ZN(n_1292));
   AND2_X1 i_1573 (.A1(b_mantissa[3]), .A2(a_mantissa[20]), .ZN(n_1295));
   INV_X1 i_1574 (.A(n_1321), .ZN(n_1299));
   NAND2_X1 i_1575 (.A1(b_mantissa[2]), .A2(a_mantissa[19]), .ZN(n_1321));
   NAND2_X1 i_1576 (.A1(b_mantissa[19]), .A2(a_mantissa[3]), .ZN(n_1325));
   AOI22_X1 i_1577 (.A1(b_mantissa[17]), .A2(a_mantissa[5]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[4]), .ZN(n_1326));
   INV_X1 i_1578 (.A(n_1329), .ZN(n_1327));
   NAND3_X1 i_1579 (.A1(b_mantissa[17]), .A2(a_mantissa[4]), .A3(n_1333), 
      .ZN(n_1329));
   AND2_X1 i_1580 (.A1(b_mantissa[18]), .A2(a_mantissa[5]), .ZN(n_1333));
   NAND2_X1 i_1581 (.A1(b_mantissa[16]), .A2(a_mantissa[6]), .ZN(n_1334));
   AOI22_X1 i_1582 (.A1(b_mantissa[14]), .A2(a_mantissa[8]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[7]), .ZN(n_1342));
   INV_X1 i_1583 (.A(n_1360), .ZN(n_1350));
   NAND3_X1 i_1584 (.A1(b_mantissa[14]), .A2(a_mantissa[7]), .A3(n_1364), 
      .ZN(n_1360));
   AND2_X1 i_1585 (.A1(b_mantissa[15]), .A2(a_mantissa[8]), .ZN(n_1364));
   NAND2_X1 i_1586 (.A1(b_mantissa[13]), .A2(a_mantissa[9]), .ZN(n_1366));
   AOI22_X1 i_1587 (.A1(b_mantissa[11]), .A2(a_mantissa[11]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[10]), .ZN(n_1374));
   NAND2_X1 i_1588 (.A1(n_1402), .A2(n_1380), .ZN(n_1376));
   AND2_X1 i_1589 (.A1(b_mantissa[12]), .A2(a_mantissa[11]), .ZN(n_1380));
   AND2_X1 i_1590 (.A1(b_mantissa[11]), .A2(a_mantissa[10]), .ZN(n_1402));
   INV_X1 i_1591 (.A(a_mantissa[1]), .ZN(n_1403));
   INV_X1 i_1592 (.A(a_mantissa[2]), .ZN(n_1407));
   INV_X1 i_1593 (.A(b_mantissa[19]), .ZN(n_1409));
   INV_X1 i_1594 (.A(b_mantissa[20]), .ZN(n_1410));
   INV_X1 i_1595 (.A(b_mantissa[21]), .ZN(n_1414));
   XNOR2_X1 i_1596 (.A(n_1427), .B(n_1424), .ZN(n_1416));
   AOI21_X1 i_1597 (.A(n_1428), .B1(n_1333), .B2(n_1430), .ZN(n_1424));
   NAND2_X1 i_1598 (.A1(a_mantissa[4]), .A2(b_mantissa[20]), .ZN(n_1427));
   AOI22_X1 i_1599 (.A1(a_mantissa[6]), .A2(b_mantissa[18]), .B1(a_mantissa[5]), 
      .B2(b_mantissa[19]), .ZN(n_1428));
   NAND2_X1 i_1600 (.A1(n_1333), .A2(n_1430), .ZN(n_1429));
   NOR2_X1 i_1601 (.A1(n_1431), .A2(n_1409), .ZN(n_1430));
   INV_X1 i_1602 (.A(a_mantissa[6]), .ZN(n_1431));
   FA_X1 i_1603 (.A(n_1531), .B(n_1524), .CI(n_1517), .CO(n_1630), .S(n_1434));
   FA_X1 i_1604 (.A(n_1630), .B(n_1624), .CI(n_1702), .CO(n_1714), .S(n_1435));
   FA_X1 i_1605 (.A(n_1603), .B(n_1596), .CI(n_1589), .CO(n_1710), .S(n_1436));
   FA_X1 i_1606 (.A(b_mantissa[2]), .B(n_1617), .CI(n_1610), .CO(n_1708), 
      .S(n_1707));
   FA_X1 i_1607 (.A(n_1659), .B(n_1710), .CI(n_1708), .CO(n_1437), .S(n_1790));
   FA_X1 i_1608 (.A(n_1602), .B(n_1595), .CI(n_1588), .CO(n_1638), .S(n_1438));
   FA_X1 i_1609 (.A(n_1623), .B(n_1616), .CI(n_1609), .CO(n_1636), .S(n_1441));
   FA_X1 i_1610 (.A(n_1707), .B(n_1638), .CI(n_1636), .CO(n_1722), .S(n_1442));
   FA_X1 i_1611 (.A(n_1714), .B(n_1790), .CI(n_1722), .CO(n_1444), .S(n_1443));
   INV_X1 i_1612 (.A(b_mantissa[7]), .ZN(n_1445));
   INV_X1 i_1613 (.A(a_mantissa[18]), .ZN(n_1448));
   NOR2_X1 i_1614 (.A1(n_1445), .A2(n_1448), .ZN(n_1449));
   NAND2_X1 i_1615 (.A1(n_1449), .A2(n_1276), .ZN(n_1450));
   INV_X1 i_1616 (.A(n_1450), .ZN(n_1451));
   AOI22_X1 i_1617 (.A1(a_mantissa[17]), .A2(b_mantissa[7]), .B1(b_mantissa[6]), 
      .B2(a_mantissa[18]), .ZN(n_1454));
   NOR2_X1 i_1618 (.A1(n_1451), .A2(n_1454), .ZN(n_1455));
   NAND2_X1 i_1619 (.A1(a_mantissa[16]), .A2(b_mantissa[8]), .ZN(n_1456));
   XNOR2_X1 i_1620 (.A(n_1455), .B(n_1456), .ZN(n_1609));
   AND2_X1 i_1621 (.A1(a_mantissa[21]), .A2(b_mantissa[4]), .ZN(n_1457));
   NAND2_X1 i_1622 (.A1(n_1457), .A2(n_1295), .ZN(n_1458));
   INV_X1 i_1623 (.A(n_1458), .ZN(n_1462));
   AOI22_X1 i_1624 (.A1(a_mantissa[20]), .A2(b_mantissa[4]), .B1(b_mantissa[3]), 
      .B2(a_mantissa[21]), .ZN(n_1466));
   NOR2_X1 i_1625 (.A1(n_1462), .A2(n_1466), .ZN(n_1468));
   NAND2_X1 i_1626 (.A1(a_mantissa[19]), .A2(b_mantissa[5]), .ZN(n_1470));
   XNOR2_X1 i_1627 (.A(n_1468), .B(n_1470), .ZN(n_1616));
   INV_X1 i_1628 (.A(b_mantissa[1]), .ZN(n_1475));
   AOI21_X1 i_1629 (.A(b_mantissa[0]), .B1(b_mantissa[1]), .B2(a_mantissa[22]), 
      .ZN(n_1476));
   AND2_X1 i_1630 (.A1(b_mantissa[0]), .A2(a_mantissa[22]), .ZN(n_1485));
   INV_X1 i_1631 (.A(n_1476), .ZN(n_1488));
   AND2_X1 i_1632 (.A1(b_mantissa[2]), .A2(a_mantissa[21]), .ZN(n_1489));
   OAI211_X1 i_1633 (.A(n_1488), .B(b_mantissa[1]), .C1(n_1489), .C2(n_1485), 
      .ZN(n_1490));
   AOI21_X1 i_1634 (.A(b_mantissa[1]), .B1(n_1489), .B2(b_mantissa[0]), .ZN(
      n_1491));
   INV_X1 i_1635 (.A(n_1491), .ZN(n_1492));
   NAND2_X1 i_1636 (.A1(n_1490), .A2(n_1492), .ZN(n_1493));
   NAND2_X1 i_1637 (.A1(b_mantissa[2]), .A2(a_mantissa[22]), .ZN(n_1494));
   XOR2_X1 i_1638 (.A(n_1493), .B(n_1494), .Z(n_1623));
   AND2_X1 i_1639 (.A1(b_mantissa[16]), .A2(a_mantissa[9]), .ZN(n_1497));
   NAND2_X1 i_1640 (.A1(n_1497), .A2(n_1364), .ZN(n_1498));
   INV_X1 i_1641 (.A(n_1498), .ZN(n_1499));
   AOI22_X1 i_1642 (.A1(a_mantissa[8]), .A2(b_mantissa[16]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[9]), .ZN(n_1500));
   NOR2_X1 i_1643 (.A1(n_1499), .A2(n_1500), .ZN(n_1501));
   NAND2_X1 i_1644 (.A1(b_mantissa[17]), .A2(a_mantissa[7]), .ZN(n_1504));
   XNOR2_X1 i_1645 (.A(n_1501), .B(n_1504), .ZN(n_1588));
   INV_X1 i_1646 (.A(b_mantissa[13]), .ZN(n_1506));
   INV_X1 i_1647 (.A(a_mantissa[12]), .ZN(n_1507));
   NOR2_X1 i_1648 (.A1(n_1506), .A2(n_1507), .ZN(n_1508));
   NAND2_X1 i_1649 (.A1(n_1508), .A2(n_1380), .ZN(n_1511));
   INV_X1 i_1650 (.A(n_1511), .ZN(n_1512));
   AOI22_X1 i_1651 (.A1(a_mantissa[11]), .A2(b_mantissa[13]), .B1(b_mantissa[12]), 
      .B2(a_mantissa[12]), .ZN(n_1513));
   NOR2_X1 i_1652 (.A1(n_1512), .A2(n_1513), .ZN(n_1514));
   NAND2_X1 i_1653 (.A1(b_mantissa[14]), .A2(a_mantissa[10]), .ZN(n_1515));
   XNOR2_X1 i_1654 (.A(n_1514), .B(n_1515), .ZN(n_1595));
   INV_X1 i_1655 (.A(a_mantissa[15]), .ZN(n_1518));
   NOR2_X1 i_1656 (.A1(n_1518), .A2(n_554), .ZN(n_1519));
   NAND2_X1 i_1657 (.A1(n_1519), .A2(n_1269), .ZN(n_1521));
   INV_X1 i_1658 (.A(n_1521), .ZN(n_1525));
   AOI22_X1 i_1659 (.A1(a_mantissa[14]), .A2(b_mantissa[10]), .B1(b_mantissa[9]), 
      .B2(a_mantissa[15]), .ZN(n_1526));
   NOR2_X1 i_1660 (.A1(n_1525), .A2(n_1526), .ZN(n_1534));
   NAND2_X1 i_1661 (.A1(a_mantissa[13]), .A2(b_mantissa[11]), .ZN(n_1541));
   XNOR2_X1 i_1662 (.A(n_1534), .B(n_1541), .ZN(n_1602));
   OAI21_X1 i_1663 (.A(n_1450), .B1(n_1454), .B2(n_1456), .ZN(n_1610));
   OAI21_X1 i_1664 (.A(n_1458), .B1(n_1466), .B2(n_1470), .ZN(n_1617));
   OAI21_X1 i_1665 (.A(n_1498), .B1(n_1500), .B2(n_1504), .ZN(n_1589));
   OAI21_X1 i_1666 (.A(n_1511), .B1(n_1513), .B2(n_1515), .ZN(n_1596));
   OAI21_X1 i_1667 (.A(n_1521), .B1(n_1526), .B2(n_1541), .ZN(n_1603));
   AOI21_X1 i_1668 (.A(a_mantissa[2]), .B1(b_mantissa[21]), .B2(a_mantissa[4]), 
      .ZN(n_1577));
   NAND3_X1 i_1669 (.A1(b_mantissa[21]), .A2(a_mantissa[2]), .A3(a_mantissa[4]), 
      .ZN(n_1578));
   NAND2_X1 i_1670 (.A1(b_mantissa[22]), .A2(a_mantissa[3]), .ZN(n_1580));
   AOI21_X1 i_1671 (.A(n_1577), .B1(n_1578), .B2(n_1580), .ZN(n_1659));
   AND2_X1 i_1672 (.A1(a_mantissa[20]), .A2(b_mantissa[5]), .ZN(n_1581));
   AND2_X1 i_1673 (.A1(a_mantissa[22]), .A2(b_mantissa[3]), .ZN(n_1583));
   NAND3_X1 i_1674 (.A1(n_1583), .A2(a_mantissa[21]), .A3(b_mantissa[4]), 
      .ZN(n_1584));
   OR2_X1 i_1675 (.A1(n_1457), .A2(n_1583), .ZN(n_1585));
   NAND2_X1 i_1676 (.A1(n_1584), .A2(n_1585), .ZN(n_1587));
   XNOR2_X1 i_1677 (.A(n_1587), .B(n_1581), .ZN(n_1702));
   AOI21_X1 i_1678 (.A(n_1491), .B1(n_1490), .B2(n_1494), .ZN(n_1624));
   NAND3_X1 i_1679 (.A1(n_1269), .A2(b_mantissa[10]), .A3(a_mantissa[13]), 
      .ZN(n_1591));
   AOI21_X1 i_1680 (.A(n_1269), .B1(b_mantissa[10]), .B2(a_mantissa[13]), 
      .ZN(n_1592));
   NAND2_X1 i_1681 (.A1(b_mantissa[11]), .A2(a_mantissa[12]), .ZN(n_1594));
   OAI21_X1 i_1682 (.A(n_1591), .B1(n_1592), .B2(n_1594), .ZN(n_1517));
   NAND3_X1 i_1683 (.A1(n_1276), .A2(b_mantissa[7]), .A3(a_mantissa[16]), 
      .ZN(n_1598));
   AOI21_X1 i_1684 (.A(n_1276), .B1(b_mantissa[7]), .B2(a_mantissa[16]), 
      .ZN(n_1599));
   NAND2_X1 i_1685 (.A1(b_mantissa[8]), .A2(a_mantissa[15]), .ZN(n_1601));
   OAI21_X1 i_1686 (.A(n_1598), .B1(n_1599), .B2(n_1601), .ZN(n_1524));
   NAND3_X1 i_1687 (.A1(n_1295), .A2(b_mantissa[4]), .A3(a_mantissa[19]), 
      .ZN(n_1605));
   AOI21_X1 i_1688 (.A(n_1295), .B1(b_mantissa[4]), .B2(a_mantissa[19]), 
      .ZN(n_1606));
   NAND2_X1 i_1689 (.A1(b_mantissa[5]), .A2(a_mantissa[18]), .ZN(n_1608));
   OAI21_X1 i_1690 (.A(n_1605), .B1(n_1606), .B2(n_1608), .ZN(n_1531));
   FA_X1 i_1691 (.A(n_1829), .B(n_1822), .CI(n_1813), .CO(n_1613), .S(n_1612));
   XNOR2_X1 i_1692 (.A(n_1619), .B(n_1614), .ZN(n_1813));
   AOI21_X1 i_1693 (.A(n_1621), .B1(a_mantissa[4]), .B2(n_1622), .ZN(n_1614));
   XNOR2_X1 i_1694 (.A(n_1625), .B(n_1615), .ZN(n_1822));
   AOI21_X1 i_1695 (.A(n_1626), .B1(n_1635), .B2(n_1628), .ZN(n_1615));
   XNOR2_X1 i_1696 (.A(n_1637), .B(n_1618), .ZN(n_1829));
   AOI21_X1 i_1697 (.A(n_1657), .B1(n_1663), .B2(n_1661), .ZN(n_1618));
   NAND2_X1 i_1698 (.A1(b_mantissa[22]), .A2(a_mantissa[5]), .ZN(n_1619));
   NAND2_X1 i_1699 (.A1(a_mantissa[4]), .A2(n_1622), .ZN(n_1620));
   NOR2_X1 i_1700 (.A1(a_mantissa[4]), .A2(n_1622), .ZN(n_1621));
   AND2_X1 i_1701 (.A1(b_mantissa[21]), .A2(a_mantissa[6]), .ZN(n_1622));
   NAND2_X1 i_1702 (.A1(b_mantissa[20]), .A2(a_mantissa[7]), .ZN(n_1625));
   AOI22_X1 i_1703 (.A1(b_mantissa[19]), .A2(a_mantissa[8]), .B1(b_mantissa[18]), 
      .B2(a_mantissa[9]), .ZN(n_1626));
   NAND2_X1 i_1704 (.A1(n_1635), .A2(n_1628), .ZN(n_1627));
   INV_X1 i_1705 (.A(n_1629), .ZN(n_1628));
   NAND2_X1 i_1706 (.A1(b_mantissa[19]), .A2(a_mantissa[9]), .ZN(n_1629));
   AND2_X1 i_1707 (.A1(b_mantissa[18]), .A2(a_mantissa[8]), .ZN(n_1635));
   NAND2_X1 i_1708 (.A1(b_mantissa[17]), .A2(a_mantissa[10]), .ZN(n_1637));
   AOI22_X1 i_1709 (.A1(b_mantissa[16]), .A2(a_mantissa[11]), .B1(b_mantissa[15]), 
      .B2(a_mantissa[12]), .ZN(n_1657));
   NAND2_X1 i_1710 (.A1(n_1663), .A2(n_1661), .ZN(n_1660));
   INV_X1 i_1711 (.A(n_1662), .ZN(n_1661));
   NAND2_X1 i_1712 (.A1(b_mantissa[16]), .A2(a_mantissa[12]), .ZN(n_1662));
   AND2_X1 i_1713 (.A1(b_mantissa[15]), .A2(a_mantissa[11]), .ZN(n_1663));
   FA_X1 i_1714 (.A(n_1905), .B(n_1898), .CI(n_1889), .CO(n_1664), .S(n_2000));
   FA_X1 i_1715 (.A(n_1926), .B(n_1919), .CI(n_1912), .CO(n_1665), .S(n_1998));
   FA_X1 i_1716 (.A(n_1911), .B(n_1904), .CI(n_1897), .CO(n_1939), .S(n_1666));
   FA_X1 i_1717 (.A(n_2000), .B(n_1998), .CI(n_1939), .CO(n_1670), .S(n_1669));
   XNOR2_X1 i_1718 (.A(n_1680), .B(n_1671), .ZN(n_1897));
   AOI21_X1 i_1719 (.A(n_1683), .B1(n_1628), .B2(n_1754), .ZN(n_1671));
   XNOR2_X1 i_1720 (.A(n_1686), .B(n_1672), .ZN(n_1904));
   AOI21_X1 i_1721 (.A(n_1687), .B1(n_1661), .B2(n_1756), .ZN(n_1672));
   XNOR2_X1 i_1722 (.A(n_1676), .B(n_1673), .ZN(n_1911));
   AOI21_X1 i_1723 (.A(n_1677), .B1(n_1704), .B2(n_1691), .ZN(n_1673));
   OAI22_X1 i_1724 (.A1(n_1706), .A2(n_1700), .B1(n_1677), .B2(n_1676), .ZN(
      n_1912));
   NAND2_X1 i_1725 (.A1(b_mantissa[14]), .A2(a_mantissa[14]), .ZN(n_1676));
   NOR2_X1 i_1726 (.A1(n_1704), .A2(n_1691), .ZN(n_1677));
   OAI21_X1 i_1727 (.A(n_1721), .B1(n_1713), .B2(n_1709), .ZN(n_1919));
   INV_X1 i_1728 (.A(n_1678), .ZN(n_1926));
   OAI21_X1 i_1729 (.A(n_1679), .B1(n_1743), .B2(n_1740), .ZN(n_1678));
   OAI21_X1 i_1730 (.A(n_1738), .B1(n_1744), .B2(n_1742), .ZN(n_1679));
   AOI21_X1 i_1731 (.A(n_1751), .B1(n_1750), .B2(n_1748), .ZN(n_1889));
   OAI21_X1 i_1732 (.A(n_1684), .B1(n_1683), .B2(n_1680), .ZN(n_1898));
   NAND2_X1 i_1733 (.A1(b_mantissa[20]), .A2(a_mantissa[8]), .ZN(n_1680));
   NOR2_X1 i_1734 (.A1(n_1757), .A2(n_1754), .ZN(n_1683));
   NAND2_X1 i_1735 (.A1(n_1628), .A2(n_1754), .ZN(n_1684));
   OAI21_X1 i_1736 (.A(n_1690), .B1(n_1687), .B2(n_1686), .ZN(n_1905));
   NAND2_X1 i_1737 (.A1(b_mantissa[17]), .A2(a_mantissa[11]), .ZN(n_1686));
   NOR2_X1 i_1738 (.A1(n_1758), .A2(n_1756), .ZN(n_1687));
   NAND2_X1 i_1739 (.A1(n_1661), .A2(n_1756), .ZN(n_1690));
   INV_X1 i_1740 (.A(n_1700), .ZN(n_1691));
   NAND2_X1 i_1741 (.A1(b_mantissa[12]), .A2(a_mantissa[16]), .ZN(n_1700));
   INV_X1 i_1742 (.A(n_1706), .ZN(n_1704));
   NAND2_X1 i_1743 (.A1(b_mantissa[13]), .A2(a_mantissa[15]), .ZN(n_1706));
   NAND2_X1 i_1744 (.A1(b_mantissa[11]), .A2(a_mantissa[17]), .ZN(n_1709));
   AOI21_X1 i_1745 (.A(n_1735), .B1(b_mantissa[10]), .B2(a_mantissa[18]), 
      .ZN(n_1713));
   NAND3_X1 i_1746 (.A1(b_mantissa[10]), .A2(a_mantissa[18]), .A3(n_1735), 
      .ZN(n_1721));
   AND2_X1 i_1747 (.A1(b_mantissa[9]), .A2(a_mantissa[19]), .ZN(n_1735));
   NAND2_X1 i_1748 (.A1(b_mantissa[8]), .A2(a_mantissa[20]), .ZN(n_1738));
   INV_X1 i_1749 (.A(n_1742), .ZN(n_1740));
   NAND2_X1 i_1750 (.A1(b_mantissa[6]), .A2(a_mantissa[22]), .ZN(n_1742));
   INV_X1 i_1751 (.A(n_1744), .ZN(n_1743));
   NAND2_X1 i_1752 (.A1(b_mantissa[7]), .A2(a_mantissa[21]), .ZN(n_1744));
   NAND2_X1 i_1753 (.A1(b_mantissa[22]), .A2(a_mantissa[6]), .ZN(n_1748));
   NAND3_X1 i_1754 (.A1(b_mantissa[21]), .A2(a_mantissa[7]), .A3(a_mantissa[5]), 
      .ZN(n_1750));
   AOI21_X1 i_1755 (.A(a_mantissa[5]), .B1(b_mantissa[21]), .B2(a_mantissa[7]), 
      .ZN(n_1751));
   AND2_X1 i_1756 (.A1(b_mantissa[18]), .A2(a_mantissa[10]), .ZN(n_1754));
   AND2_X1 i_1757 (.A1(b_mantissa[15]), .A2(a_mantissa[13]), .ZN(n_1756));
   INV_X1 i_1758 (.A(n_1629), .ZN(n_1757));
   INV_X1 i_1759 (.A(n_1662), .ZN(n_1758));
   FA_X1 i_1760 (.A(n_271), .B(n_270), .CI(n_269), .CO(n_268), .S(n_1761));
   FA_X1 i_1761 (.A(n_274), .B(n_272), .CI(n_268), .CO(n_1764), .S(n_1763));
   OAI22_X1 i_1762 (.A1(n_957), .A2(n_1770), .B1(n_1768), .B2(n_1765), .ZN(n_269));
   OAI21_X1 i_1763 (.A(n_1785), .B1(n_1784), .B2(n_1772), .ZN(n_270));
   AOI22_X1 i_1764 (.A1(n_1818), .A2(n_1816), .B1(n_1800), .B2(n_1791), .ZN(
      n_271));
   AOI21_X1 i_1765 (.A(n_1824), .B1(n_1821), .B2(n_1819), .ZN(n_272));
   AOI21_X1 i_1766 (.A(n_1828), .B1(n_1832), .B2(n_1827), .ZN(n_274));
   NAND2_X1 i_1767 (.A1(b_mantissa[22]), .A2(a_mantissa[15]), .ZN(n_1765));
   AOI21_X1 i_1768 (.A(a_mantissa[14]), .B1(b_mantissa[21]), .B2(a_mantissa[16]), 
      .ZN(n_1768));
   NAND2_X1 i_1769 (.A1(b_mantissa[21]), .A2(a_mantissa[14]), .ZN(n_1770));
   NAND2_X1 i_1770 (.A1(b_mantissa[20]), .A2(a_mantissa[17]), .ZN(n_1772));
   AOI22_X1 i_1771 (.A1(b_mantissa[18]), .A2(a_mantissa[19]), .B1(b_mantissa[19]), 
      .B2(a_mantissa[18]), .ZN(n_1784));
   NAND4_X1 i_1772 (.A1(b_mantissa[18]), .A2(a_mantissa[19]), .A3(b_mantissa[19]), 
      .A4(a_mantissa[18]), .ZN(n_1785));
   NAND2_X1 i_1773 (.A1(b_mantissa[17]), .A2(a_mantissa[20]), .ZN(n_1791));
   INV_X1 i_1774 (.A(n_1801), .ZN(n_1800));
   NOR2_X1 i_1775 (.A1(n_1818), .A2(n_1816), .ZN(n_1801));
   NAND2_X1 i_1776 (.A1(b_mantissa[15]), .A2(a_mantissa[22]), .ZN(n_1816));
   NAND2_X1 i_1777 (.A1(b_mantissa[16]), .A2(a_mantissa[21]), .ZN(n_1818));
   NAND2_X1 i_1778 (.A1(b_mantissa[22]), .A2(a_mantissa[16]), .ZN(n_1819));
   NAND3_X1 i_1779 (.A1(b_mantissa[21]), .A2(a_mantissa[17]), .A3(a_mantissa[15]), 
      .ZN(n_1821));
   AOI21_X1 i_1780 (.A(a_mantissa[15]), .B1(b_mantissa[21]), .B2(a_mantissa[17]), 
      .ZN(n_1824));
   NAND2_X1 i_1781 (.A1(b_mantissa[20]), .A2(a_mantissa[18]), .ZN(n_1827));
   INV_X1 i_1782 (.A(n_1831), .ZN(n_1828));
   OAI21_X1 i_1783 (.A(n_1835), .B1(n_1409), .B2(n_1198), .ZN(n_1831));
   NAND4_X1 i_1784 (.A1(b_mantissa[18]), .A2(a_mantissa[20]), .A3(b_mantissa[19]), 
      .A4(a_mantissa[19]), .ZN(n_1832));
   NAND2_X1 i_1785 (.A1(b_mantissa[18]), .A2(a_mantissa[20]), .ZN(n_1835));
   FA_X1 i_1786 (.A(n_302), .B(n_285), .CI(n_275), .CO(n_1839), .S(n_1838));
   XNOR2_X1 i_1787 (.A(n_1900), .B(n_1871), .ZN(n_275));
   OAI22_X1 i_1788 (.A1(n_1198), .A2(n_1901), .B1(a_mantissa[19]), .B2(n_1938), 
      .ZN(n_1871));
   XNOR2_X1 i_1789 (.A(n_1999), .B(n_1872), .ZN(n_285));
   NOR2_X1 i_1790 (.A1(n_2009), .A2(n_2001), .ZN(n_1872));
   AOI22_X1 i_1791 (.A1(n_2105), .A2(n_1894), .B1(n_1448), .B2(n_2110), .ZN(
      n_302));
   NAND2_X1 i_1792 (.A1(a_mantissa[18]), .A2(n_2107), .ZN(n_1894));
   NAND2_X1 i_1793 (.A1(b_mantissa[22]), .A2(a_mantissa[20]), .ZN(n_1900));
   INV_X1 i_1794 (.A(n_1938), .ZN(n_1901));
   NAND2_X1 i_1795 (.A1(b_mantissa[21]), .A2(a_mantissa[21]), .ZN(n_1938));
   NAND2_X1 i_1796 (.A1(b_mantissa[20]), .A2(a_mantissa[22]), .ZN(n_1999));
   AOI21_X1 i_1797 (.A(b_mantissa[19]), .B1(b_mantissa[18]), .B2(n_2097), 
      .ZN(n_2001));
   INV_X1 i_1798 (.A(n_2009), .ZN(n_2008));
   AOI211_X1 i_1799 (.A(n_1409), .B(n_2104), .C1(n_2099), .C2(n_2098), .ZN(
      n_2009));
   INV_X1 i_1800 (.A(n_2098), .ZN(n_2097));
   NAND2_X1 i_1801 (.A1(b_mantissa[20]), .A2(a_mantissa[21]), .ZN(n_2098));
   NAND2_X1 i_1802 (.A1(b_mantissa[18]), .A2(a_mantissa[22]), .ZN(n_2099));
   INV_X1 i_1803 (.A(n_2104), .ZN(n_2103));
   AOI21_X1 i_1804 (.A(b_mantissa[18]), .B1(b_mantissa[19]), .B2(a_mantissa[22]), 
      .ZN(n_2104));
   NAND2_X1 i_1805 (.A1(b_mantissa[22]), .A2(a_mantissa[19]), .ZN(n_2105));
   INV_X1 i_1806 (.A(n_2110), .ZN(n_2107));
   NAND2_X1 i_1807 (.A1(b_mantissa[21]), .A2(a_mantissa[20]), .ZN(n_2110));
endmodule

module datapath__0_3(p_0, p_1, O_final_mantessa);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]O_final_mantessa;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(O_final_mantessa[0]));
   HA_X1 i_1 (.A(p_1[1]), .B(n_0), .CO(n_1), .S(O_final_mantessa[1]));
   HA_X1 i_2 (.A(p_1[2]), .B(n_1), .CO(n_2), .S(O_final_mantessa[2]));
   HA_X1 i_3 (.A(p_1[3]), .B(n_2), .CO(n_3), .S(O_final_mantessa[3]));
   HA_X1 i_4 (.A(p_1[4]), .B(n_3), .CO(n_4), .S(O_final_mantessa[4]));
   HA_X1 i_5 (.A(p_1[5]), .B(n_4), .CO(n_5), .S(O_final_mantessa[5]));
   HA_X1 i_6 (.A(p_1[6]), .B(n_5), .CO(n_6), .S(O_final_mantessa[6]));
   HA_X1 i_7 (.A(p_1[7]), .B(n_6), .CO(n_7), .S(O_final_mantessa[7]));
   HA_X1 i_8 (.A(p_1[8]), .B(n_7), .CO(n_8), .S(O_final_mantessa[8]));
   HA_X1 i_9 (.A(p_1[9]), .B(n_8), .CO(n_9), .S(O_final_mantessa[9]));
   HA_X1 i_10 (.A(p_1[10]), .B(n_9), .CO(n_10), .S(O_final_mantessa[10]));
   HA_X1 i_11 (.A(p_1[11]), .B(n_10), .CO(n_11), .S(O_final_mantessa[11]));
   HA_X1 i_12 (.A(p_1[12]), .B(n_11), .CO(n_12), .S(O_final_mantessa[12]));
   HA_X1 i_13 (.A(p_1[13]), .B(n_12), .CO(n_13), .S(O_final_mantessa[13]));
   HA_X1 i_14 (.A(p_1[14]), .B(n_13), .CO(n_14), .S(O_final_mantessa[14]));
   HA_X1 i_15 (.A(p_1[15]), .B(n_14), .CO(n_15), .S(O_final_mantessa[15]));
   HA_X1 i_16 (.A(p_1[16]), .B(n_15), .CO(n_16), .S(O_final_mantessa[16]));
   HA_X1 i_17 (.A(p_1[17]), .B(n_16), .CO(n_17), .S(O_final_mantessa[17]));
   HA_X1 i_18 (.A(p_1[18]), .B(n_17), .CO(n_18), .S(O_final_mantessa[18]));
   HA_X1 i_19 (.A(p_1[19]), .B(n_18), .CO(n_19), .S(O_final_mantessa[19]));
   HA_X1 i_20 (.A(p_1[20]), .B(n_19), .CO(n_20), .S(O_final_mantessa[20]));
   HA_X1 i_21 (.A(p_1[21]), .B(n_20), .CO(n_21), .S(O_final_mantessa[21]));
   XOR2_X1 i_22 (.A(p_1[22]), .B(n_21), .Z(O_final_mantessa[22]));
endmodule

module FloatingPointMultiplier(A, B, O, OF);
   input [31:0]A;
   input [31:0]B;
   output [31:0]O;
   output OF;

   wire [47:0]o_mantissa;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_1_15;
   wire n_0_1_16;
   wire n_0_1_24;
   wire n_0_1_17;
   wire n_0_1_25;
   wire n_0_1_18;
   wire n_0_1_26;
   wire n_0_1_19;
   wire n_0_1_27;
   wire n_0_1_20;
   wire n_0_1_28;
   wire n_0_1_21;
   wire n_0_1_29;
   wire n_0_1_22;
   wire n_0_1_30;
   wire n_0_1_23;
   wire n_0_1_14;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_34;
   wire n_0_1_35;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_1_103;
   wire n_0_1_104;
   wire n_0_1_31;
   wire n_0_1_32;
   wire n_0_1_33;
   wire n_0_1_36;
   wire n_0_1_37;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_1_60;
   wire n_0_1_61;
   wire n_0_1_62;
   wire n_0_1_63;
   wire n_0_1_64;
   wire n_0_23;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_105;

   datapath i_0_0 (.b_mantissa({1'b1, B[22], B[21], B[20], B[19], B[18], B[17], 
      B[16], B[15], B[14], B[13], B[12], B[11], B[10], B[9], B[8], B[7], B[6], 
      B[5], B[4], B[3], B[2], B[1], B[0]}), .a_mantissa({1'b1, A[22], A[21], 
      A[20], A[19], A[18], A[17], A[16], A[15], A[14], A[13], A[12], A[11], 
      A[10], A[9], A[8], A[7], A[6], A[5], A[4], A[3], A[2], A[1], A[0]}), 
      .o_mantissa(o_mantissa));
   datapath__0_3 i_0_5 (.p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, n_0_23}), .p_1({n_0_46, n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, 
      n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, 
      n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24}), 
      .O_final_mantessa({n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0}));
   HA_X1 i_0_1_0 (.A(B[24]), .B(A[24]), .CO(n_0_1_3), .S(n_0_1_2));
   HA_X1 i_0_1_1 (.A(B[25]), .B(A[25]), .CO(n_0_1_5), .S(n_0_1_4));
   HA_X1 i_0_1_2 (.A(B[26]), .B(A[26]), .CO(n_0_1_7), .S(n_0_1_6));
   HA_X1 i_0_1_3 (.A(B[27]), .B(A[27]), .CO(n_0_1_9), .S(n_0_1_8));
   HA_X1 i_0_1_4 (.A(B[28]), .B(A[28]), .CO(n_0_1_11), .S(n_0_1_10));
   HA_X1 i_0_1_5 (.A(B[29]), .B(A[29]), .CO(n_0_1_13), .S(n_0_1_12));
   HA_X1 i_0_1_6 (.A(A[23]), .B(n_0_1_0), .CO(n_0_1_16), .S(n_0_1_15));
   FA_X1 i_0_1_7 (.A(n_0_1_1), .B(n_0_1_2), .CI(n_0_1_16), .CO(n_0_1_17), 
      .S(n_0_1_24));
   FA_X1 i_0_1_8 (.A(n_0_1_3), .B(n_0_1_4), .CI(n_0_1_17), .CO(n_0_1_18), 
      .S(n_0_1_25));
   FA_X1 i_0_1_9 (.A(n_0_1_5), .B(n_0_1_6), .CI(n_0_1_18), .CO(n_0_1_19), 
      .S(n_0_1_26));
   FA_X1 i_0_1_10 (.A(n_0_1_7), .B(n_0_1_8), .CI(n_0_1_19), .CO(n_0_1_20), 
      .S(n_0_1_27));
   FA_X1 i_0_1_11 (.A(n_0_1_9), .B(n_0_1_10), .CI(n_0_1_20), .CO(n_0_1_21), 
      .S(n_0_1_28));
   FA_X1 i_0_1_12 (.A(n_0_1_11), .B(n_0_1_12), .CI(n_0_1_21), .CO(n_0_1_22), 
      .S(n_0_1_29));
   FA_X1 i_0_1_13 (.A(n_0_1_13), .B(n_0_1_14), .CI(n_0_1_22), .CO(n_0_1_23), 
      .S(n_0_1_30));
   XNOR2_X1 i_0_1_14 (.A(B[30]), .B(A[30]), .ZN(n_0_1_14));
   XNOR2_X1 i_0_1_15 (.A(B[23]), .B(o_mantissa[47]), .ZN(n_0_1_0));
   OR2_X1 i_0_1_16 (.A1(B[23]), .A2(o_mantissa[47]), .ZN(n_0_1_1));
   OAI21_X1 i_0_1_17 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_82), .ZN(O[0]));
   OAI21_X1 i_0_1_21 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_83), .ZN(O[1]));
   OAI21_X1 i_0_1_22 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_84), .ZN(O[2]));
   OAI21_X1 i_0_1_23 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_85), .ZN(O[3]));
   OAI21_X1 i_0_1_24 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_86), .ZN(O[4]));
   OAI21_X1 i_0_1_25 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_87), .ZN(O[5]));
   OAI21_X1 i_0_1_26 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_88), .ZN(O[6]));
   OAI21_X1 i_0_1_27 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_89), .ZN(O[7]));
   OAI21_X1 i_0_1_28 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_90), .ZN(O[8]));
   OAI21_X1 i_0_1_29 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_91), .ZN(O[9]));
   OAI21_X1 i_0_1_30 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_92), .ZN(O[10]));
   OAI21_X1 i_0_1_31 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_93), .ZN(O[11]));
   OAI21_X1 i_0_1_32 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_94), .ZN(O[12]));
   OAI21_X1 i_0_1_33 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_95), .ZN(O[13]));
   OAI21_X1 i_0_1_34 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_96), .ZN(O[14]));
   OAI21_X1 i_0_1_35 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_97), .ZN(O[15]));
   OAI21_X1 i_0_1_36 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_98), .ZN(O[16]));
   OAI21_X1 i_0_1_37 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_99), .ZN(O[17]));
   OAI21_X1 i_0_1_38 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_100), .ZN(O[18]));
   OAI21_X1 i_0_1_39 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_101), .ZN(O[19]));
   OAI21_X1 i_0_1_40 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_102), .ZN(O[20]));
   OAI21_X1 i_0_1_41 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_103), .ZN(O[21]));
   OAI21_X1 i_0_1_42 (.A(n_0_1_34), .B1(n_0_1_33), .B2(n_0_1_104), .ZN(O[22]));
   AOI221_X1 i_0_1_18 (.A(n_0_1_35), .B1(n_0_1_42), .B2(n_0_1_59), .C1(n_0_1_62), 
      .C2(n_0_1_50), .ZN(n_0_1_34));
   NOR2_X1 i_0_1_19 (.A1(n_0_1_58), .A2(n_0_1_36), .ZN(n_0_1_35));
   OAI21_X1 i_0_1_20 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_81), .ZN(O[23]));
   OAI21_X1 i_0_1_47 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_80), .ZN(O[24]));
   OAI21_X1 i_0_1_48 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_79), .ZN(O[25]));
   OAI21_X1 i_0_1_49 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_78), .ZN(O[26]));
   OAI21_X1 i_0_1_50 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_77), .ZN(O[27]));
   OAI21_X1 i_0_1_51 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_76), .ZN(O[28]));
   OAI21_X1 i_0_1_52 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_75), .ZN(O[29]));
   OAI21_X1 i_0_1_53 (.A(n_0_1_58), .B1(n_0_1_37), .B2(n_0_1_74), .ZN(O[30]));
   XOR2_X1 i_0_1_83 (.A(B[31]), .B(A[31]), .Z(O[31]));
   MUX2_X1 i_0_1_94 (.A(o_mantissa[23]), .B(o_mantissa[24]), .S(o_mantissa[47]), 
      .Z(n_0_24));
   MUX2_X1 i_0_1_95 (.A(o_mantissa[24]), .B(o_mantissa[25]), .S(o_mantissa[47]), 
      .Z(n_0_25));
   MUX2_X1 i_0_1_96 (.A(o_mantissa[25]), .B(o_mantissa[26]), .S(o_mantissa[47]), 
      .Z(n_0_26));
   MUX2_X1 i_0_1_97 (.A(o_mantissa[26]), .B(o_mantissa[27]), .S(o_mantissa[47]), 
      .Z(n_0_27));
   MUX2_X1 i_0_1_98 (.A(o_mantissa[27]), .B(o_mantissa[28]), .S(o_mantissa[47]), 
      .Z(n_0_28));
   MUX2_X1 i_0_1_99 (.A(o_mantissa[28]), .B(o_mantissa[29]), .S(o_mantissa[47]), 
      .Z(n_0_29));
   MUX2_X1 i_0_1_100 (.A(o_mantissa[29]), .B(o_mantissa[30]), .S(o_mantissa[47]), 
      .Z(n_0_30));
   MUX2_X1 i_0_1_101 (.A(o_mantissa[30]), .B(o_mantissa[31]), .S(o_mantissa[47]), 
      .Z(n_0_31));
   MUX2_X1 i_0_1_102 (.A(o_mantissa[31]), .B(o_mantissa[32]), .S(o_mantissa[47]), 
      .Z(n_0_32));
   MUX2_X1 i_0_1_103 (.A(o_mantissa[32]), .B(o_mantissa[33]), .S(o_mantissa[47]), 
      .Z(n_0_33));
   MUX2_X1 i_0_1_104 (.A(o_mantissa[33]), .B(o_mantissa[34]), .S(o_mantissa[47]), 
      .Z(n_0_34));
   MUX2_X1 i_0_1_105 (.A(o_mantissa[34]), .B(o_mantissa[35]), .S(o_mantissa[47]), 
      .Z(n_0_35));
   MUX2_X1 i_0_1_106 (.A(o_mantissa[35]), .B(o_mantissa[36]), .S(o_mantissa[47]), 
      .Z(n_0_36));
   MUX2_X1 i_0_1_107 (.A(o_mantissa[36]), .B(o_mantissa[37]), .S(o_mantissa[47]), 
      .Z(n_0_37));
   MUX2_X1 i_0_1_108 (.A(o_mantissa[37]), .B(o_mantissa[38]), .S(o_mantissa[47]), 
      .Z(n_0_38));
   MUX2_X1 i_0_1_109 (.A(o_mantissa[38]), .B(o_mantissa[39]), .S(o_mantissa[47]), 
      .Z(n_0_39));
   MUX2_X1 i_0_1_110 (.A(o_mantissa[39]), .B(o_mantissa[40]), .S(o_mantissa[47]), 
      .Z(n_0_40));
   MUX2_X1 i_0_1_111 (.A(o_mantissa[40]), .B(o_mantissa[41]), .S(o_mantissa[47]), 
      .Z(n_0_41));
   MUX2_X1 i_0_1_112 (.A(o_mantissa[41]), .B(o_mantissa[42]), .S(o_mantissa[47]), 
      .Z(n_0_42));
   MUX2_X1 i_0_1_113 (.A(o_mantissa[42]), .B(o_mantissa[43]), .S(o_mantissa[47]), 
      .Z(n_0_43));
   MUX2_X1 i_0_1_114 (.A(o_mantissa[43]), .B(o_mantissa[44]), .S(o_mantissa[47]), 
      .Z(n_0_44));
   MUX2_X1 i_0_1_115 (.A(o_mantissa[44]), .B(o_mantissa[45]), .S(o_mantissa[47]), 
      .Z(n_0_45));
   MUX2_X1 i_0_1_116 (.A(o_mantissa[45]), .B(o_mantissa[46]), .S(o_mantissa[47]), 
      .Z(n_0_46));
   INV_X1 i_0_1_117 (.A(n_0_1_30), .ZN(n_0_1_74));
   INV_X1 i_0_1_118 (.A(n_0_1_29), .ZN(n_0_1_75));
   INV_X1 i_0_1_119 (.A(n_0_1_28), .ZN(n_0_1_76));
   INV_X1 i_0_1_120 (.A(n_0_1_27), .ZN(n_0_1_77));
   INV_X1 i_0_1_121 (.A(n_0_1_26), .ZN(n_0_1_78));
   INV_X1 i_0_1_122 (.A(n_0_1_25), .ZN(n_0_1_79));
   INV_X1 i_0_1_123 (.A(n_0_1_24), .ZN(n_0_1_80));
   INV_X1 i_0_1_43 (.A(n_0_1_15), .ZN(n_0_1_81));
   INV_X1 i_0_1_44 (.A(n_0_0), .ZN(n_0_1_82));
   INV_X1 i_0_1_126 (.A(n_0_1), .ZN(n_0_1_83));
   INV_X1 i_0_1_127 (.A(n_0_2), .ZN(n_0_1_84));
   INV_X1 i_0_1_128 (.A(n_0_3), .ZN(n_0_1_85));
   INV_X1 i_0_1_129 (.A(n_0_4), .ZN(n_0_1_86));
   INV_X1 i_0_1_130 (.A(n_0_5), .ZN(n_0_1_87));
   INV_X1 i_0_1_131 (.A(n_0_6), .ZN(n_0_1_88));
   INV_X1 i_0_1_132 (.A(n_0_7), .ZN(n_0_1_89));
   INV_X1 i_0_1_133 (.A(n_0_8), .ZN(n_0_1_90));
   INV_X1 i_0_1_134 (.A(n_0_9), .ZN(n_0_1_91));
   INV_X1 i_0_1_135 (.A(n_0_10), .ZN(n_0_1_92));
   INV_X1 i_0_1_136 (.A(n_0_11), .ZN(n_0_1_93));
   INV_X1 i_0_1_137 (.A(n_0_12), .ZN(n_0_1_94));
   INV_X1 i_0_1_138 (.A(n_0_13), .ZN(n_0_1_95));
   INV_X1 i_0_1_139 (.A(n_0_14), .ZN(n_0_1_96));
   INV_X1 i_0_1_140 (.A(n_0_15), .ZN(n_0_1_97));
   INV_X1 i_0_1_141 (.A(n_0_16), .ZN(n_0_1_98));
   INV_X1 i_0_1_142 (.A(n_0_17), .ZN(n_0_1_99));
   INV_X1 i_0_1_143 (.A(n_0_18), .ZN(n_0_1_100));
   INV_X1 i_0_1_144 (.A(n_0_19), .ZN(n_0_1_101));
   INV_X1 i_0_1_145 (.A(n_0_20), .ZN(n_0_1_102));
   INV_X1 i_0_1_146 (.A(n_0_21), .ZN(n_0_1_103));
   INV_X1 i_0_1_147 (.A(n_0_22), .ZN(n_0_1_104));
   AOI211_X1 i_0_1_45 (.A(n_0_1_31), .B(n_0_1_33), .C1(n_0_1_23), .C2(n_0_1_32), 
      .ZN(OF));
   NOR2_X1 i_0_1_46 (.A1(n_0_1_23), .A2(n_0_1_32), .ZN(n_0_1_31));
   NOR2_X1 i_0_1_54 (.A1(A[30]), .A2(B[30]), .ZN(n_0_1_32));
   NAND2_X1 i_0_1_55 (.A1(n_0_1_58), .A2(n_0_1_36), .ZN(n_0_1_33));
   INV_X1 i_0_1_56 (.A(n_0_1_37), .ZN(n_0_1_36));
   OAI33_X1 i_0_1_57 (.A1(n_0_1_41), .A2(n_0_1_40), .A3(n_0_1_42), .B1(n_0_1_39), 
      .B2(n_0_1_38), .B3(n_0_1_50), .ZN(n_0_1_37));
   OR4_X1 i_0_1_58 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(n_0_1_38));
   OR4_X1 i_0_1_59 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(n_0_1_39));
   OR4_X1 i_0_1_60 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(n_0_1_40));
   OR4_X1 i_0_1_61 (.A1(B[25]), .A2(B[24]), .A3(B[26]), .A4(B[23]), .ZN(n_0_1_41));
   NAND3_X1 i_0_1_62 (.A1(n_0_1_49), .A2(n_0_1_48), .A3(n_0_1_43), .ZN(n_0_1_42));
   AND4_X1 i_0_1_63 (.A1(n_0_1_47), .A2(n_0_1_46), .A3(n_0_1_45), .A4(n_0_1_44), 
      .ZN(n_0_1_43));
   NOR4_X1 i_0_1_64 (.A1(B[6]), .A2(B[5]), .A3(B[4]), .A4(B[3]), .ZN(n_0_1_44));
   NOR3_X1 i_0_1_65 (.A1(B[2]), .A2(B[1]), .A3(B[0]), .ZN(n_0_1_45));
   NOR4_X1 i_0_1_66 (.A1(B[14]), .A2(B[13]), .A3(B[12]), .A4(B[11]), .ZN(
      n_0_1_46));
   NOR4_X1 i_0_1_67 (.A1(B[10]), .A2(B[9]), .A3(B[8]), .A4(B[7]), .ZN(n_0_1_47));
   NOR4_X1 i_0_1_68 (.A1(B[22]), .A2(B[19]), .A3(B[17]), .A4(B[16]), .ZN(
      n_0_1_48));
   NOR4_X1 i_0_1_69 (.A1(B[21]), .A2(B[20]), .A3(B[18]), .A4(B[15]), .ZN(
      n_0_1_49));
   NAND3_X1 i_0_1_70 (.A1(n_0_1_57), .A2(n_0_1_56), .A3(n_0_1_51), .ZN(n_0_1_50));
   AND4_X1 i_0_1_71 (.A1(n_0_1_55), .A2(n_0_1_54), .A3(n_0_1_53), .A4(n_0_1_52), 
      .ZN(n_0_1_51));
   NOR4_X1 i_0_1_72 (.A1(A[6]), .A2(A[5]), .A3(A[4]), .A4(A[3]), .ZN(n_0_1_52));
   NOR3_X1 i_0_1_73 (.A1(A[2]), .A2(A[1]), .A3(A[0]), .ZN(n_0_1_53));
   NOR4_X1 i_0_1_74 (.A1(A[14]), .A2(A[13]), .A3(A[12]), .A4(A[11]), .ZN(
      n_0_1_54));
   NOR4_X1 i_0_1_75 (.A1(A[10]), .A2(A[9]), .A3(A[8]), .A4(A[7]), .ZN(n_0_1_55));
   NOR4_X1 i_0_1_76 (.A1(A[22]), .A2(A[19]), .A3(A[17]), .A4(A[16]), .ZN(
      n_0_1_56));
   NOR4_X1 i_0_1_77 (.A1(A[21]), .A2(A[20]), .A3(A[18]), .A4(A[15]), .ZN(
      n_0_1_57));
   NOR2_X1 i_0_1_78 (.A1(n_0_1_62), .A2(n_0_1_59), .ZN(n_0_1_58));
   NOR2_X1 i_0_1_79 (.A1(n_0_1_61), .A2(n_0_1_60), .ZN(n_0_1_59));
   NAND4_X1 i_0_1_80 (.A1(B[30]), .A2(B[29]), .A3(B[28]), .A4(B[27]), .ZN(
      n_0_1_60));
   NAND4_X1 i_0_1_81 (.A1(B[26]), .A2(B[25]), .A3(B[24]), .A4(B[23]), .ZN(
      n_0_1_61));
   NOR2_X1 i_0_1_82 (.A1(n_0_1_64), .A2(n_0_1_63), .ZN(n_0_1_62));
   NAND4_X1 i_0_1_84 (.A1(A[30]), .A2(A[29]), .A3(A[28]), .A4(A[27]), .ZN(
      n_0_1_63));
   NAND4_X1 i_0_1_85 (.A1(A[26]), .A2(A[25]), .A3(A[24]), .A4(A[23]), .ZN(
      n_0_1_64));
   INV_X1 i_0_1_86 (.A(n_0_1_65), .ZN(n_0_23));
   OAI222_X1 i_0_1_87 (.A1(n_0_1_105), .A2(o_mantissa[23]), .B1(o_mantissa[47]), 
      .B2(o_mantissa[22]), .C1(n_0_1_71), .C2(n_0_1_66), .ZN(n_0_1_65));
   NAND4_X1 i_0_1_88 (.A1(n_0_1_70), .A2(n_0_1_69), .A3(n_0_1_68), .A4(n_0_1_67), 
      .ZN(n_0_1_66));
   NOR4_X1 i_0_1_89 (.A1(o_mantissa[6]), .A2(o_mantissa[5]), .A3(o_mantissa[4]), 
      .A4(o_mantissa[3]), .ZN(n_0_1_67));
   NOR3_X1 i_0_1_90 (.A1(o_mantissa[2]), .A2(o_mantissa[1]), .A3(o_mantissa[0]), 
      .ZN(n_0_1_68));
   NOR4_X1 i_0_1_91 (.A1(o_mantissa[14]), .A2(o_mantissa[13]), .A3(
      o_mantissa[12]), .A4(o_mantissa[11]), .ZN(n_0_1_69));
   NOR4_X1 i_0_1_92 (.A1(o_mantissa[10]), .A2(o_mantissa[9]), .A3(o_mantissa[8]), 
      .A4(o_mantissa[7]), .ZN(n_0_1_70));
   NAND2_X1 i_0_1_93 (.A1(n_0_1_73), .A2(n_0_1_72), .ZN(n_0_1_71));
   NOR4_X1 i_0_1_124 (.A1(o_mantissa[22]), .A2(o_mantissa[19]), .A3(
      o_mantissa[17]), .A4(o_mantissa[16]), .ZN(n_0_1_72));
   NOR4_X1 i_0_1_125 (.A1(o_mantissa[21]), .A2(o_mantissa[20]), .A3(
      o_mantissa[18]), .A4(o_mantissa[15]), .ZN(n_0_1_73));
   INV_X1 i_0_1_148 (.A(o_mantissa[47]), .ZN(n_0_1_105));
endmodule
