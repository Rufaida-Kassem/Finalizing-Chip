* SPICE NETLIST
***************************************

.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT WELLTAP
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_2
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT ICV_3
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=3 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKGATETST_X1 SE E CK VDD VSS GCK 7
** N=19 EP=7 IP=0 FDC=24
M0 8 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=205 $D=1
M1 VSS E 8 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.94e-14 PD=8.3e-07 PS=7e-07 $X=335 $Y=205 $D=1
M2 17 8 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=525 $Y=140 $D=1
M3 9 12 17 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.915e-14 AS=3.85e-14 PD=9.1e-07 PS=8.3e-07 $X=715 $Y=140 $D=1
M4 18 10 9 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.915e-14 PD=4.6e-07 PS=9.1e-07 $X=945 $Y=300 $D=1
M5 VSS 11 18 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=1135 $Y=300 $D=1
M6 10 12 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=1325 $Y=180 $D=1
M7 VSS 9 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1665 $Y=315 $D=1
M8 12 CK VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1855 $Y=315 $D=1
M9 19 CK 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=2240 $Y=295 $D=1
M10 VSS 9 19 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.835e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2430 $Y=295 $D=1
M11 GCK 13 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.835e-14 PD=6e-07 PS=7e-07 $X=2620 $Y=310 $D=1
M12 14 SE 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=890 $D=0
M13 VDD E 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=4.41e-14 PD=1.12e-06 PS=9.1e-07 $X=335 $Y=890 $D=0
M14 15 8 VDD VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=525 $Y=890 $D=0
M15 9 10 15 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=3.93e-14 AS=5.88e-14 PD=1.2e-06 PS=1.12e-06 $X=715 $Y=890 $D=0
M16 16 12 9 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.93e-14 PD=4.6e-07 PS=1.2e-06 $X=945 $Y=990 $D=0
M17 VDD 11 16 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=1135 $Y=990 $D=0
M18 10 12 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=1325 $Y=990 $D=0
M19 VDD 9 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1665 $Y=870 $D=0
M20 12 CK VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1855 $Y=870 $D=0
M21 13 CK VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=2240 $Y=870 $D=0
M22 VDD 9 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2430 $Y=870 $D=0
M23 GCK 13 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2620 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN
** N=7 EP=5 IP=0 FDC=6
M0 6 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 6 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 6 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT ICV_7
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q
** N=20 EP=5 IP=0 FDC=28
M0 VSS 9 6 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 17 8 VSS VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 7 6 17 VSS NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 18 9 7 VSS NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 18 VSS NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 8 7 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 19 7 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 10 6 19 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 20 9 10 VSS NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 12 20 VSS NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 12 10 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 10 QN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 12 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 9 6 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 13 8 VDD VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 7 9 13 VDD PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 14 6 7 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 14 VDD PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 8 7 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 15 7 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 10 9 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 16 6 10 VDD PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 12 16 VDD PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 12 10 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 10 QN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 12 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_8
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6
** N=8 EP=6 IP=0 FDC=6
M0 8 A1 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 7 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD
** N=8 EP=6 IP=0 FDC=6
M0 ZN B2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 7 B1 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 8 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=2 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5
** N=5 EP=5 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=3 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7
** N=13 EP=7 IP=0 FDC=16
M0 12 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 12 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 9 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 9 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 13 A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 10 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 8 A S VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 9 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 9 A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 10 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 10 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT INV_X2 A ZN VSS VDD
** N=4 EP=4 IP=0 FDC=4
M0 ZN A VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6
** N=10 EP=6 IP=0 FDC=10
M0 7 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 10 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 10 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 9 A 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 8 B Z VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 42 43 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95
** N=179 EP=93 IP=2357 FDC=1400
X1057 35 117 32 34 35 17 35 CLKGATETST_X1 $T=72630 82200 1 0 $X=72515 $Y=80685
X1058 35 118 32 34 35 26 35 CLKGATETST_X1 $T=74150 85000 1 0 $X=74035 $Y=83485
X1059 35 121 32 34 35 1 35 CLKGATETST_X1 $T=81560 82200 0 0 $X=81445 $Y=82085
X1116 63 31 35 34 117 OR2_X1 $T=73200 82200 1 180 $X=72325 $Y=82085
X1117 63 31 35 34 118 OR2_X1 $T=73390 85000 1 0 $X=73275 $Y=83485
X1118 63 31 35 34 121 OR2_X1 $T=80230 85000 1 0 $X=80115 $Y=83485
X1170 78 1 35 34 74 DFF_X1 $T=5560 79400 1 180 $X=2215 $Y=79285
X1171 157 1 35 34 65 DFF_X1 $T=5560 82200 0 180 $X=2215 $Y=80685
X1172 142 1 35 34 36 DFF_X1 $T=2330 85000 1 0 $X=2215 $Y=83485
X1173 158 1 35 34 37 DFF_X1 $T=5560 85000 1 0 $X=5445 $Y=83485
X1174 174 1 35 34 79 DFF_X1 $T=10310 82200 0 180 $X=6965 $Y=80685
X1175 170 1 35 34 38 DFF_X1 $T=8790 85000 1 0 $X=8675 $Y=83485
X1176 171 1 35 34 80 DFF_X1 $T=14300 82200 1 0 $X=14185 $Y=80685
X1177 172 1 35 34 81 DFF_X1 $T=15440 85000 1 0 $X=15325 $Y=83485
X1178 122 1 35 34 39 DFF_X1 $T=18290 82200 1 0 $X=18175 $Y=80685
X1179 159 1 35 34 66 DFF_X1 $T=18670 85000 1 0 $X=18555 $Y=83485
X1180 160 1 35 34 82 DFF_X1 $T=22280 85000 1 0 $X=22165 $Y=83485
X1181 161 1 35 34 76 DFF_X1 $T=25510 85000 1 0 $X=25395 $Y=83485
X1182 105 1 35 34 56 DFF_X1 $T=28740 85000 1 0 $X=28625 $Y=83485
X1183 107 1 35 34 43 DFF_X1 $T=31970 85000 1 0 $X=31855 $Y=83485
X1184 162 17 35 34 34 DFF_X1 $T=36720 79400 0 0 $X=36605 $Y=79285
X1185 109 1 35 34 83 DFF_X1 $T=37860 85000 1 0 $X=37745 $Y=83485
X1186 133 26 35 34 57 DFF_X1 $T=38620 82200 1 0 $X=38505 $Y=80685
X1187 123 26 35 34 58 DFF_X1 $T=43750 82200 1 0 $X=43635 $Y=80685
X1188 164 26 35 34 59 DFF_X1 $T=45460 85000 1 0 $X=45345 $Y=83485
X1189 163 26 35 34 71 DFF_X1 $T=46980 82200 1 0 $X=46865 $Y=80685
X1190 135 1 35 34 84 DFF_X1 $T=48690 85000 1 0 $X=48575 $Y=83485
X1191 137 1 35 34 72 DFF_X1 $T=55530 85000 1 0 $X=55415 $Y=83485
X1192 151 1 35 34 85 DFF_X1 $T=58760 85000 1 0 $X=58645 $Y=83485
X1193 140 1 35 34 49 DFF_X1 $T=62370 85000 1 0 $X=62255 $Y=83485
X1194 167 1 35 34 86 DFF_X1 $T=70160 85000 1 0 $X=70045 $Y=83485
X1195 173 1 35 34 62 DFF_X1 $T=77000 85000 1 0 $X=76885 $Y=83485
X1196 169 1 35 34 64 DFF_X1 $T=78710 79400 0 0 $X=78595 $Y=79285
X1197 168 1 35 34 73 DFF_X1 $T=78710 82200 1 0 $X=78595 $Y=80685
X1218 12 2 35 34 142 35 AND2_X1 $T=5370 82200 0 0 $X=5255 $Y=82085
X1219 12 97 35 34 157 35 AND2_X1 $T=6320 82200 0 180 $X=5445 $Y=80685
X1220 12 98 35 34 158 35 AND2_X1 $T=7080 82200 0 180 $X=6205 $Y=80685
X1221 12 99 35 34 174 35 AND2_X1 $T=9550 79400 1 180 $X=8675 $Y=79285
X1222 12 4 35 34 170 35 AND2_X1 $T=11070 79400 0 0 $X=10955 $Y=79285
X1223 12 5 35 34 171 35 AND2_X1 $T=14110 79400 1 180 $X=13235 $Y=79285
X1224 12 100 35 34 172 35 AND2_X1 $T=15250 79400 0 0 $X=15135 $Y=79285
X1225 12 101 35 34 159 35 AND2_X1 $T=17530 82200 1 0 $X=17415 $Y=80685
X1226 12 6 35 34 122 35 AND2_X1 $T=20190 79400 1 180 $X=19315 $Y=79285
X1227 12 102 35 34 160 35 AND2_X1 $T=23420 82200 0 180 $X=22545 $Y=80685
X1228 12 103 35 34 161 35 AND2_X1 $T=25510 82200 1 0 $X=25395 $Y=80685
X1229 33 9 35 34 40 35 AND2_X1 $T=27790 82200 1 0 $X=27675 $Y=80685
X1230 12 104 35 34 105 35 AND2_X1 $T=28740 82200 0 0 $X=28625 $Y=82085
X1231 45 10 35 34 55 35 AND2_X1 $T=29500 82200 1 0 $X=29385 $Y=80685
X1232 12 106 35 34 107 35 AND2_X1 $T=31400 82200 1 0 $X=31285 $Y=80685
X1233 12 108 35 34 109 35 AND2_X1 $T=34060 82200 1 0 $X=33945 $Y=80685
X1234 33 14 35 34 42 35 AND2_X1 $T=35390 79400 1 180 $X=34515 $Y=79285
X1235 33 15 35 34 68 35 AND2_X1 $T=35580 82200 1 0 $X=35465 $Y=80685
X1236 33 16 35 34 162 35 AND2_X1 $T=36340 82200 1 0 $X=36225 $Y=80685
X1237 45 18 35 34 133 35 AND2_X1 $T=38620 82200 0 0 $X=38505 $Y=82085
X1238 45 20 35 34 69 35 AND2_X1 $T=41090 82200 0 0 $X=40975 $Y=82085
X1239 45 21 35 34 77 35 AND2_X1 $T=41090 85000 1 0 $X=40975 $Y=83485
X1240 45 22 35 34 47 35 AND2_X1 $T=42990 82200 0 180 $X=42115 $Y=80685
X1241 45 46 35 34 70 35 AND2_X1 $T=42990 82200 1 0 $X=42875 $Y=80685
X1242 45 23 35 34 123 35 AND2_X1 $T=42990 85000 1 0 $X=42875 $Y=83485
X1243 45 24 35 34 163 35 AND2_X1 $T=44700 82200 0 0 $X=44585 $Y=82085
X1244 45 25 35 34 164 35 AND2_X1 $T=44700 85000 1 0 $X=44585 $Y=83485
X1245 12 110 35 34 135 35 AND2_X1 $T=51160 82200 1 180 $X=50285 $Y=82085
X1246 12 111 35 34 137 35 AND2_X1 $T=54770 82200 0 0 $X=54655 $Y=82085
X1247 12 112 35 34 151 35 AND2_X1 $T=58570 82200 0 0 $X=58455 $Y=82085
X1248 12 113 35 34 140 35 AND2_X1 $T=62370 82200 0 0 $X=62255 $Y=82085
X1249 12 114 35 34 167 35 AND2_X1 $T=66550 82200 1 0 $X=66435 $Y=80685
X1250 12 115 35 34 168 35 AND2_X1 $T=69780 82200 1 0 $X=69665 $Y=80685
X1251 12 116 35 34 173 35 AND2_X1 $T=69970 82200 0 0 $X=69855 $Y=82085
X1252 12 119 35 34 61 35 AND2_X1 $T=75480 79400 0 0 $X=75365 $Y=79285
X1253 12 120 35 34 169 35 AND2_X1 $T=75480 82200 1 0 $X=75365 $Y=80685
X1351 50 3 98 51 35 34 OAI21_X1 $T=6890 79400 0 0 $X=6775 $Y=79285
X1352 126 3 97 51 35 34 OAI21_X1 $T=8410 79400 1 180 $X=7535 $Y=79285
X1353 127 3 99 51 35 34 OAI21_X1 $T=10310 79400 1 180 $X=9435 $Y=79285
X1354 87 3 100 51 35 34 OAI21_X1 $T=16010 79400 0 0 $X=15895 $Y=79285
X1355 128 3 101 51 35 34 OAI21_X1 $T=18100 79400 1 180 $X=17225 $Y=79285
X1356 143 7 102 53 35 34 OAI21_X1 $T=23420 82200 1 0 $X=23305 $Y=80685
X1357 175 7 103 53 35 34 OAI21_X1 $T=25320 82200 0 0 $X=25205 $Y=82085
X1358 129 7 104 53 35 34 OAI21_X1 $T=27790 82200 0 180 $X=26915 $Y=80685
X1359 146 7 106 53 35 34 OAI21_X1 $T=30640 82200 1 0 $X=30525 $Y=80685
X1360 132 7 108 53 35 34 OAI21_X1 $T=34060 82200 0 180 $X=33185 $Y=80685
X1361 124 7 110 53 35 34 OAI21_X1 $T=47740 82200 0 0 $X=47625 $Y=82085
X1362 165 7 111 53 35 34 OAI21_X1 $T=53060 82200 0 0 $X=52945 $Y=82085
X1363 125 7 112 53 35 34 OAI21_X1 $T=56670 82200 0 0 $X=56555 $Y=82085
X1364 177 7 113 53 35 34 OAI21_X1 $T=61230 82200 0 0 $X=61115 $Y=82085
X1365 153 7 114 53 35 34 OAI21_X1 $T=65410 82200 1 0 $X=65295 $Y=80685
X1366 154 7 115 53 35 34 OAI21_X1 $T=67310 82200 1 0 $X=67195 $Y=80685
X1367 166 7 116 53 35 34 OAI21_X1 $T=68830 82200 0 180 $X=67955 $Y=80685
X1368 155 7 120 53 35 34 OAI21_X1 $T=71300 82200 0 180 $X=70425 $Y=80685
X1369 141 7 119 53 35 34 OAI21_X1 $T=73960 79400 0 0 $X=73845 $Y=79285
X1392 88 35 34 126 35 INV_X1 $T=8790 79400 1 180 $X=8295 $Y=79285
X1393 89 35 34 127 35 INV_X1 $T=11070 79400 1 180 $X=10575 $Y=79285
X1394 90 35 34 128 35 INV_X1 $T=18480 79400 1 180 $X=17985 $Y=79285
X1395 91 35 34 143 35 INV_X1 $T=23420 79400 0 0 $X=23305 $Y=79285
X1396 67 35 34 175 35 INV_X1 $T=25130 82200 1 0 $X=25015 $Y=80685
X1397 144 35 34 129 35 INV_X1 $T=26650 82200 1 0 $X=26535 $Y=80685
X1398 145 35 34 146 35 INV_X1 $T=30260 82200 1 0 $X=30145 $Y=80685
X1399 147 35 34 132 35 INV_X1 $T=32920 82200 1 0 $X=32805 $Y=80685
X1400 31 35 34 33 35 INV_X1 $T=41850 82200 0 0 $X=41735 $Y=82085
X1401 134 35 34 124 35 INV_X1 $T=45840 82200 0 0 $X=45725 $Y=82085
X1402 148 35 34 165 35 INV_X1 $T=52490 82200 1 0 $X=52375 $Y=80685
X1403 149 35 34 125 35 INV_X1 $T=55720 82200 1 0 $X=55605 $Y=80685
X1404 150 35 34 177 35 INV_X1 $T=58760 82200 1 0 $X=58645 $Y=80685
X1405 152 35 34 153 35 INV_X1 $T=63510 82200 1 0 $X=63395 $Y=80685
X1406 31 35 34 12 35 INV_X1 $T=64840 82200 0 0 $X=64725 $Y=82085
X1407 179 35 34 166 35 INV_X1 $T=66170 82200 1 0 $X=66055 $Y=80685
X1408 48 35 34 154 35 INV_X1 $T=66360 79400 0 0 $X=66245 $Y=79285
X1409 92 35 34 155 35 INV_X1 $T=69210 79400 0 0 $X=69095 $Y=79285
X1410 93 35 34 141 35 INV_X1 $T=72060 79400 0 0 $X=71945 $Y=79285
X1473 144 176 8 35 34 54 35 HA_X1 $T=27030 79400 0 0 $X=26915 $Y=79285
X1474 145 130 11 35 34 176 35 HA_X1 $T=30830 79400 1 180 $X=28815 $Y=79285
X1475 147 131 13 35 34 130 35 HA_X1 $T=32730 79400 1 180 $X=30715 $Y=79285
X1476 134 156 19 35 34 131 35 HA_X1 $T=39950 79400 0 0 $X=39835 $Y=79285
X1477 148 136 27 35 34 156 35 HA_X1 $T=53440 79400 0 0 $X=53325 $Y=79285
X1478 149 138 28 35 34 136 35 HA_X1 $T=57240 79400 1 180 $X=55225 $Y=79285
X1479 150 139 29 35 34 138 35 HA_X1 $T=59140 79400 1 180 $X=57125 $Y=79285
X1480 152 178 94 35 34 139 35 HA_X1 $T=59900 82200 1 0 $X=59785 $Y=80685
X1481 179 60 30 35 34 178 35 HA_X1 $T=64270 79400 1 180 $X=62255 $Y=79285
X1492 31 45 35 34 INV_X2 $T=44320 85000 0 180 $X=43635 $Y=83485
X1510 34 75 52 95 35 35 XOR2_X1 $T=23420 79400 1 180 $X=22165 $Y=79285
.ENDS
***************************************
.SUBCKT MUX2_X1 A S B VSS VDD Z
** N=12 EP=6 IP=0 FDC=12
M0 VSS S 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 11 A VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 8 7 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 12 S 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=715 $Y=90 $D=1
M4 VSS B 12 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=905 $Y=90 $D=1
M5 Z 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 VDD S 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M7 9 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M8 8 S 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M9 10 7 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=715 $Y=995 $D=0
M10 VDD B 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=905 $Y=995 $D=0
M11 Z 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6
** N=7 EP=6 IP=0 FDC=4
M0 7 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 7 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6
** N=7 EP=6 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 7 A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 7 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD 7
** N=9 EP=7 IP=0 FDC=6
M0 9 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 8 B1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN 7
** N=9 EP=7 IP=0 FDC=6
M0 ZN A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 9 A2 8 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6
** N=10 EP=6 IP=0 FDC=10
M0 10 A 7 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 10 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 8 7 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 8 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 7 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 9 A ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN
** N=9 EP=6 IP=0 FDC=8
M0 VSS A1 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 7 A2 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 7 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 7 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 8 A1 7 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 9 A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 7 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD
** N=10 EP=7 IP=0 FDC=8
M0 VSS B2 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 8 B1 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 8 A2 ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 10 A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS 8
** N=11 EP=8 IP=0 FDC=8
M0 ZN A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 9 A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 10 A3 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 11 A2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 11 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8
** N=20 EP=8 IP=0 FDC=28
M0 VSS 9 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 18 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 9 A 18 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 10 CI 9 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 10 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 12 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 12 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 14 9 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 19 CI 14 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 20 B 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 14 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 9 CO VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 15 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 9 A 15 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 11 CI 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 11 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 13 B VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 13 A VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 14 9 13 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 16 CI 14 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 17 B 16 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 17 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 14 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143
** N=256 EP=143 IP=2758 FDC=1508
X1294 72 6 34 33 251 OR2_X1 $T=20380 76600 1 180 $X=19505 $Y=76485
X1326 113 1 34 33 194 DFF_X1 $T=1000 73800 0 0 $X=885 $Y=73685
X1327 34 11 34 33 245 DFF_X1 $T=2330 76600 0 0 $X=2215 $Y=76485
X1328 114 11 34 33 58 DFF_X1 $T=26650 73800 0 0 $X=26535 $Y=73685
X1329 115 1 34 33 107 DFF_X1 $T=28170 76600 1 0 $X=28055 $Y=75085
X1330 116 11 34 33 94 DFF_X1 $T=35200 76600 1 0 $X=35085 $Y=75085
X1331 117 11 34 33 60 DFF_X1 $T=35960 79400 1 0 $X=35845 $Y=77885
X1332 118 1 34 33 109 DFF_X1 $T=40520 79400 1 0 $X=40405 $Y=77885
X1333 119 1 34 33 110 DFF_X1 $T=42230 76600 1 0 $X=42115 $Y=75085
X1334 120 1 34 33 77 DFF_X1 $T=42230 76600 0 0 $X=42115 $Y=76485
X1335 18 1 34 33 111 DFF_X1 $T=43750 79400 1 0 $X=43635 $Y=77885
X1336 121 32 34 33 69 DFF_X1 $T=77950 79400 1 0 $X=77835 $Y=77885
X1337 240 32 34 33 70 DFF_X1 $T=78710 76600 0 0 $X=78595 $Y=76485
X1338 249 32 34 33 71 DFF_X1 $T=81180 73800 0 0 $X=81065 $Y=73685
X1339 217 32 34 33 112 DFF_X1 $T=81180 79400 1 0 $X=81065 $Y=77885
X1340 45 153 34 33 47 34 AND2_X1 $T=5560 79400 0 180 $X=4685 $Y=77885
X1341 38 13 34 33 92 34 AND2_X1 $T=32920 76600 0 0 $X=32805 $Y=76485
X1342 78 19 34 33 40 34 AND2_X1 $T=45460 76600 1 0 $X=45345 $Y=75085
X1343 41 166 34 33 200 34 AND2_X1 $T=47170 73800 0 0 $X=47055 $Y=73685
X1344 45 193 34 33 240 34 AND2_X1 $T=74910 76600 0 0 $X=74795 $Y=76485
X1345 45 184 34 33 104 34 AND2_X1 $T=76810 73800 1 180 $X=75935 $Y=73685
X1346 45 185 34 33 68 34 AND2_X1 $T=76810 73800 0 0 $X=76695 $Y=73685
X1347 45 186 34 33 217 34 AND2_X1 $T=77190 79400 1 0 $X=77075 $Y=77885
X1348 45 187 34 33 249 34 AND2_X1 $T=77380 76600 1 0 $X=77265 $Y=75085
X1349 45 188 34 33 105 34 AND2_X1 $T=78520 73800 0 0 $X=78405 $Y=73685
X1443 219 2 86 36 34 33 OAI21_X1 $T=6890 79400 1 0 $X=6775 $Y=77885
X1444 221 2 88 36 34 33 OAI21_X1 $T=12970 79400 1 0 $X=12855 $Y=77885
X1445 222 2 89 36 34 33 OAI21_X1 $T=14490 79400 0 180 $X=13615 $Y=77885
X1446 227 7 90 44 34 33 OAI21_X1 $T=20760 79400 0 180 $X=19885 $Y=77885
X1447 125 17 199 62 34 33 OAI21_X1 $T=41090 73800 0 0 $X=40975 $Y=73685
X1448 43 23 97 174 34 33 OAI21_X1 $T=56670 73800 0 0 $X=56555 $Y=73685
X1449 246 7 193 44 34 33 OAI21_X1 $T=65410 76600 0 0 $X=65295 $Y=76485
X1450 234 7 184 44 34 33 OAI21_X1 $T=72440 76600 1 0 $X=72325 $Y=75085
X1451 237 7 187 44 34 33 OAI21_X1 $T=74340 76600 1 0 $X=74225 $Y=75085
X1452 215 7 185 44 34 33 OAI21_X1 $T=74530 73800 0 0 $X=74415 $Y=73685
X1453 239 7 186 44 34 33 OAI21_X1 $T=75480 79400 0 180 $X=74605 $Y=77885
X1454 241 7 188 44 34 33 OAI21_X1 $T=75860 76600 0 180 $X=74985 $Y=75085
X1455 216 7 103 44 34 33 OAI21_X1 $T=76050 73800 1 180 $X=75175 $Y=73685
X1488 35 34 33 219 34 INV_X1 $T=6510 79400 1 0 $X=6395 $Y=77885
X1489 189 34 33 48 34 INV_X1 $T=8030 79400 0 180 $X=7535 $Y=77885
X1490 220 34 33 221 34 INV_X1 $T=12590 79400 1 0 $X=12475 $Y=77885
X1491 223 34 33 222 34 INV_X1 $T=14870 79400 0 180 $X=14375 $Y=77885
X1492 225 34 33 122 34 INV_X1 $T=15820 79400 1 0 $X=15705 $Y=77885
X1493 8 34 33 51 34 INV_X1 $T=20570 73800 0 0 $X=20455 $Y=73685
X1494 130 34 33 227 34 INV_X1 $T=21140 79400 0 180 $X=20645 $Y=77885
X1495 198 34 33 164 34 INV_X1 $T=37480 73800 1 180 $X=36985 $Y=73685
X1496 230 34 33 205 34 INV_X1 $T=50590 76600 0 0 $X=50475 $Y=76485
X1497 209 34 33 173 34 INV_X1 $T=55150 76600 1 180 $X=54655 $Y=76485
X1498 80 34 33 177 34 INV_X1 $T=58190 76600 1 0 $X=58075 $Y=75085
X1499 255 34 33 246 34 INV_X1 $T=60280 76600 0 0 $X=60165 $Y=76485
X1500 231 34 33 241 34 INV_X1 $T=66740 76600 1 0 $X=66625 $Y=75085
X1501 248 34 33 234 34 INV_X1 $T=67690 76600 1 0 $X=67575 $Y=75085
X1502 211 34 33 216 34 INV_X1 $T=68070 76600 1 0 $X=67955 $Y=75085
X1503 212 34 33 215 34 INV_X1 $T=72440 73800 0 0 $X=72325 $Y=73685
X1504 236 34 33 237 34 INV_X1 $T=73200 76600 1 0 $X=73085 $Y=75085
X1505 238 34 33 239 34 INV_X1 $T=74340 79400 1 0 $X=74225 $Y=77885
X1618 190 134 3 34 33 195 34 HA_X1 $T=11450 73800 1 180 $X=9435 $Y=73685
X1619 224 136 4 34 33 196 34 HA_X1 $T=15820 73800 1 180 $X=13805 $Y=73685
X1620 256 5 137 34 33 242 34 HA_X1 $T=17720 73800 1 180 $X=15705 $Y=73685
X1621 223 226 138 34 33 243 34 HA_X1 $T=19240 76600 0 180 $X=17225 $Y=75085
X1622 132 228 252 34 33 123 34 HA_X1 $T=24180 79400 0 180 $X=22165 $Y=77885
X1623 57 83 253 34 33 228 34 HA_X1 $T=26080 79400 0 180 $X=24065 $Y=77885
X1624 255 191 177 34 33 247 34 HA_X1 $T=59330 76600 1 0 $X=59215 $Y=75085
X1625 231 247 33 34 33 210 34 HA_X1 $T=61230 76600 1 0 $X=61115 $Y=75085
X1626 248 210 141 34 33 250 34 HA_X1 $T=62370 76600 0 0 $X=62255 $Y=76485
X1627 211 250 181 34 33 100 34 HA_X1 $T=63700 73800 0 0 $X=63585 $Y=73685
X1628 101 232 180 34 33 65 34 HA_X1 $T=65600 79400 0 180 $X=63585 $Y=77885
X1629 102 213 233 34 33 232 34 HA_X1 $T=67500 79400 0 180 $X=65485 $Y=77885
X1630 212 66 142 34 33 214 34 HA_X1 $T=68640 73800 0 0 $X=68525 $Y=73685
X1631 67 235 182 34 33 213 34 HA_X1 $T=71680 79400 0 180 $X=69665 $Y=77885
X1632 236 214 31 34 33 254 34 HA_X1 $T=70540 76600 1 0 $X=70425 $Y=75085
X1633 238 254 183 34 33 235 34 HA_X1 $T=73580 79400 0 180 $X=71565 $Y=77885
X1703 33 245 153 194 34 34 XOR2_X1 $T=3850 76600 1 0 $X=3735 $Y=75085
X1704 33 53 161 55 34 34 XOR2_X1 $T=26650 73800 1 180 $X=25395 $Y=73685
X1705 33 197 165 84 34 34 XOR2_X1 $T=35200 76600 0 180 $X=33945 $Y=75085
X1706 33 198 167 229 34 34 XOR2_X1 $T=39570 76600 0 180 $X=38315 $Y=75085
X1707 33 16 168 199 34 34 XOR2_X1 $T=44890 73800 0 0 $X=44775 $Y=73685
X1708 33 206 178 207 34 34 XOR2_X1 $T=54960 79400 0 180 $X=53705 $Y=77885
X1709 33 209 179 244 34 34 XOR2_X1 $T=58190 79400 1 0 $X=58075 $Y=77885
X1710 159 6 9 34 33 252 MUX2_X1 $T=23610 76600 1 180 $X=22165 $Y=76485
X1711 9 6 10 34 33 37 MUX2_X1 $T=22850 76600 1 0 $X=22735 $Y=75085
X1712 160 6 159 34 33 253 MUX2_X1 $T=23610 76600 0 0 $X=23495 $Y=76485
X1713 161 6 160 34 33 91 MUX2_X1 $T=24940 76600 0 0 $X=24825 $Y=76485
X1714 12 6 161 34 33 143 MUX2_X1 $T=28550 79400 1 0 $X=28435 $Y=77885
X1715 163 6 12 34 33 75 MUX2_X1 $T=32920 76600 1 180 $X=31475 $Y=76485
X1716 165 6 163 34 33 61 MUX2_X1 $T=39190 79400 1 0 $X=39075 $Y=77885
X1717 167 6 165 34 33 95 MUX2_X1 $T=49640 79400 0 180 $X=48195 $Y=77885
X1718 168 6 167 34 33 96 MUX2_X1 $T=49640 79400 1 0 $X=49525 $Y=77885
X1719 46 6 20 34 33 191 MUX2_X1 $T=50400 73800 0 0 $X=50285 $Y=73685
X1720 176 6 168 34 33 98 MUX2_X1 $T=58190 79400 0 180 $X=56745 $Y=77885
X1721 178 6 176 34 33 64 MUX2_X1 $T=60660 79400 0 180 $X=59215 $Y=77885
X1722 20 6 24 34 33 33 MUX2_X1 $T=60660 73800 0 0 $X=60545 $Y=73685
X1723 179 6 178 34 33 99 MUX2_X1 $T=60660 79400 1 0 $X=60545 $Y=77885
X1724 25 6 27 34 33 181 MUX2_X1 $T=62370 73800 0 0 $X=62255 $Y=73685
X1725 26 6 179 34 33 180 MUX2_X1 $T=62370 79400 1 0 $X=62255 $Y=77885
X1726 28 6 26 34 33 233 MUX2_X1 $T=67500 76600 1 180 $X=66055 $Y=76485
X1727 29 6 28 34 33 182 MUX2_X1 $T=68830 76600 0 0 $X=68715 $Y=76485
X1728 30 6 29 34 33 183 MUX2_X1 $T=70540 73800 0 0 $X=70425 $Y=73685
X1729 128 34 36 7 33 34 NAND2_X1 $T=17720 73800 0 0 $X=17605 $Y=73685
X1730 42 34 63 230 33 34 NAND2_X1 $T=51540 76600 1 180 $X=50855 $Y=76485
X1731 79 34 22 175 33 34 NAND2_X1 $T=56290 76600 0 180 $X=55605 $Y=75085
X1732 43 34 23 174 33 34 NAND2_X1 $T=58000 73800 1 180 $X=57315 $Y=73685
X1733 56 33 131 55 34 34 NOR2_X1 $T=24370 73800 1 180 $X=23685 $Y=73685
X1734 166 33 41 169 34 34 NOR2_X1 $T=47360 76600 1 0 $X=47245 $Y=75085
X1735 230 33 169 201 34 34 NOR2_X1 $T=49450 76600 1 0 $X=49335 $Y=75085
X1736 200 33 169 202 34 34 NOR2_X1 $T=49640 76600 0 0 $X=49525 $Y=76485
X1737 42 33 63 170 34 34 NOR2_X1 $T=51540 76600 1 0 $X=51425 $Y=75085
X1738 205 33 170 207 34 34 NOR2_X1 $T=52490 76600 0 0 $X=52375 $Y=76485
X1739 79 33 22 171 34 34 NOR2_X1 $T=56290 76600 1 0 $X=56175 $Y=75085
X1740 43 33 23 208 34 34 NOR2_X1 $T=56860 76600 1 0 $X=56745 $Y=75085
X1741 164 14 197 93 34 33 34 AOI21_X1 $T=34630 73800 0 0 $X=34515 $Y=73685
X1742 124 15 229 93 34 33 34 AOI21_X1 $T=37100 73800 1 180 $X=36225 $Y=73685
X1743 62 16 198 108 34 33 34 AOI21_X1 $T=38620 73800 0 0 $X=38505 $Y=73685
X1744 173 175 206 171 34 33 34 AOI21_X1 $T=54010 76600 0 0 $X=53895 $Y=76485
X1745 175 174 203 192 34 33 34 AOI21_X1 $T=54960 76600 0 180 $X=54085 $Y=75085
X1746 174 21 209 208 34 33 34 AOI21_X1 $T=54960 76600 1 0 $X=54845 $Y=75085
X1747 79 22 244 171 34 33 34 AOI21_X1 $T=57430 76600 1 180 $X=56555 $Y=76485
X1748 21 33 208 192 34 204 34 NOR3_X1 $T=54580 73800 1 180 $X=53705 $Y=73685
X1749 34 72 226 6 33 34 XNOR2_X1 $T=20380 76600 0 180 $X=19125 $Y=75085
X1750 34 129 159 158 33 34 XNOR2_X1 $T=20380 76600 1 0 $X=20265 $Y=75085
X1751 34 73 160 82 33 34 XNOR2_X1 $T=24370 73800 0 0 $X=24255 $Y=73685
X1752 34 74 163 162 33 34 XNOR2_X1 $T=31400 73800 0 0 $X=31285 $Y=73685
X1753 34 202 176 172 33 34 XNOR2_X1 $T=53820 79400 0 180 $X=52565 $Y=77885
X1754 169 170 171 34 33 192 OR3_X1 $T=52110 76600 1 0 $X=51995 $Y=75085
X1755 51 52 34 158 53 54 33 OAI22_X1 $T=20950 73800 0 0 $X=20835 $Y=73685
X1756 197 76 34 162 59 39 33 OAI22_X1 $T=32540 73800 0 0 $X=32425 $Y=73685
X1757 206 205 34 172 63 42 33 OAI22_X1 $T=52490 76600 1 180 $X=51425 $Y=76485
X1759 204 33 203 201 200 16 34 34 NOR4_X1 $T=50400 73800 1 180 $X=49335 $Y=73685
X1760 106 218 133 126 33 34 189 34 FA_X1 $T=4230 73800 0 0 $X=4115 $Y=73685
X1761 218 154 81 195 33 34 87 34 FA_X1 $T=5560 76600 0 0 $X=5445 $Y=76485
X1762 154 155 190 127 33 34 49 34 FA_X1 $T=8030 79400 1 0 $X=7915 $Y=77885
X1763 155 156 135 196 33 34 220 34 FA_X1 $T=11260 76600 1 0 $X=11145 $Y=75085
X1764 156 157 224 242 33 34 225 34 FA_X1 $T=14300 76600 1 0 $X=14185 $Y=75085
X1765 157 243 256 251 33 34 50 34 FA_X1 $T=16960 79400 1 0 $X=16845 $Y=77885
X1766 17 140 85 139 33 34 166 34 FA_X1 $T=41850 73800 0 0 $X=41735 $Y=73685
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN
** N=8 EP=6 IP=0 FDC=6
M0 7 A3 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 8 A2 7 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z
** N=5 EP=4 IP=0 FDC=4
M0 VSS A 5 VSS NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 5 VSS VSS NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 5 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 5 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN
** N=12 EP=8 IP=0 FDC=10
M0 11 B2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 11 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 12 C2 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 12 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 9 B1 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 10 A 9 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 10 VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 10 C1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 8 A1 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 8 A3 VSS VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 9 A1 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 10 A2 9 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 11 A3 10 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 11 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD
** N=10 EP=7 IP=0 FDC=8
M0 8 A4 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 9 A3 8 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 10 A2 9 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 10 VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 69 70 71 72 73 74 75 76 77 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178
** N=302 EP=175 IP=2983 FDC=1540
M0 225 223 46 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=15790 $Y=71090 $D=1
M1 46 226 225 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15980 $Y=71090 $D=1
M2 225 51 46 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16170 $Y=71090 $D=1
M3 198 18 225 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16360 $Y=71090 $D=1
M4 225 227 198 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=16550 $Y=71090 $D=1
M5 198 228 225 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=16740 $Y=71090 $D=1
M6 230 60 46 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=24895 $Y=68290 $D=1
M7 46 201 230 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=25085 $Y=68290 $D=1
M8 28 230 46 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=25275 $Y=68290 $D=1
M9 46 230 28 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=25465 $Y=68290 $D=1
M10 234 69 46 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=48845 $Y=68290 $D=1
M11 46 70 234 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=49035 $Y=68290 $D=1
M12 234 28 235 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=49400 $Y=68290 $D=1
M13 235 29 234 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=49590 $Y=68290 $D=1
M14 71 30 235 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=49780 $Y=68290 $D=1
M15 235 213 71 46 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=49970 $Y=68290 $D=1
M16 295 223 52 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=15790 $Y=71680 $D=0
M17 296 226 295 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15980 $Y=71680 $D=0
M18 198 51 296 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16170 $Y=71680 $D=0
M19 297 18 198 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16360 $Y=71680 $D=0
M20 298 227 297 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=16550 $Y=71680 $D=0
M21 52 228 298 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=16740 $Y=71680 $D=0
M22 299 60 230 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=24895 $Y=68880 $D=0
M23 52 201 299 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=25085 $Y=68880 $D=0
M24 28 230 52 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=25275 $Y=68880 $D=0
M25 52 230 28 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=25465 $Y=68880 $D=0
M26 300 69 52 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=48845 $Y=68880 $D=0
M27 71 70 300 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=49035 $Y=68880 $D=0
M28 301 28 71 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=49400 $Y=68880 $D=0
M29 52 29 301 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=49590 $Y=68880 $D=0
M30 302 30 52 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=49780 $Y=68880 $D=0
M31 71 213 302 52 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=49970 $Y=68880 $D=0
X1426 142 3 46 52 197 DFF_X1 $T=1000 68200 0 0 $X=885 $Y=68085
X1427 11 3 46 52 14 DFF_X1 $T=12400 68200 0 0 $X=12285 $Y=68085
X1428 143 44 46 52 103 DFF_X1 $T=78710 71000 1 0 $X=78595 $Y=69485
X1429 293 44 46 52 120 DFF_X1 $T=78710 71000 0 0 $X=78595 $Y=70885
X1430 144 44 46 52 121 DFF_X1 $T=78710 73800 1 0 $X=78595 $Y=72285
X1431 292 44 46 52 77 DFF_X1 $T=81180 68200 0 0 $X=81065 $Y=68085
X1452 80 1 46 52 130 46 AND2_X1 $T=1190 71000 0 0 $X=1075 $Y=70885
X1453 45 2 46 52 46 46 AND2_X1 $T=1190 73800 1 0 $X=1075 $Y=72285
X1454 20 19 46 52 229 46 AND2_X1 $T=18860 68200 0 0 $X=18745 $Y=68085
X1455 251 206 46 52 269 46 AND2_X1 $T=29310 71000 1 180 $X=28435 $Y=70885
X1456 75 222 46 52 292 46 AND2_X1 $T=77570 73800 0 180 $X=76695 $Y=72285
X1457 76 42 46 52 101 46 AND2_X1 $T=77950 68200 0 0 $X=77835 $Y=68085
X1458 75 43 46 52 293 46 AND2_X1 $T=77950 73800 1 0 $X=77835 $Y=72285
X1581 19 20 231 83 46 52 OAI21_X1 $T=19240 71000 0 0 $X=19125 $Y=70885
X1582 248 22 201 265 46 52 OAI21_X1 $T=23610 68200 1 180 $X=22735 $Y=68085
X1583 89 203 285 202 46 52 OAI21_X1 $T=26840 71000 0 180 $X=25965 $Y=69485
X1584 41 220 290 102 46 52 OAI21_X1 $T=73390 68200 1 180 $X=72515 $Y=68085
X1585 260 240 291 238 46 52 OAI21_X1 $T=73580 71000 1 180 $X=72705 $Y=70885
X1586 280 79 222 54 46 52 OAI21_X1 $T=73960 73800 1 0 $X=73845 $Y=72285
X1634 105 46 52 53 46 INV_X1 $T=18670 73800 0 180 $X=18175 $Y=72285
X1635 266 46 52 87 46 INV_X1 $T=25130 73800 0 180 $X=24635 $Y=72285
X1636 254 46 52 63 46 INV_X1 $T=32160 73800 1 0 $X=32045 $Y=72285
X1637 28 46 52 213 46 INV_X1 $T=49830 71000 1 0 $X=49715 $Y=69485
X1638 279 46 52 280 46 INV_X1 $T=69020 73800 1 0 $X=68905 $Y=72285
X1639 118 46 52 259 46 INV_X1 $T=72820 71000 0 180 $X=72325 $Y=69485
X1640 41 46 52 260 46 INV_X1 $T=75100 71000 1 0 $X=74985 $Y=69485
X1742 131 5 197 46 52 263 46 HA_X1 $T=10690 71000 1 180 $X=8675 $Y=70885
X1743 132 6 7 46 52 145 46 HA_X1 $T=11070 73800 0 180 $X=9055 $Y=72285
X1744 48 50 10 46 52 146 46 HA_X1 $T=12970 73800 0 180 $X=10955 $Y=72285
X1745 279 167 219 46 52 154 46 HA_X1 $T=65980 73800 1 0 $X=65865 $Y=72285
X1844 52 204 61 285 46 46 XOR2_X1 $T=27600 73800 1 0 $X=27485 $Y=72285
X1845 52 137 96 129 46 46 XOR2_X1 $T=56480 73800 1 0 $X=56365 $Y=72285
X1846 52 259 40 221 46 46 XOR2_X1 $T=72630 73800 0 180 $X=71375 $Y=72285
X1847 33 28 34 46 52 138 MUX2_X1 $T=60660 73800 1 0 $X=60545 $Y=72285
X1848 35 28 36 46 52 219 MUX2_X1 $T=64650 73800 1 0 $X=64535 $Y=72285
X1849 36 28 37 46 52 73 MUX2_X1 $T=67500 71000 0 0 $X=67385 $Y=70885
X1850 37 28 40 46 52 141 MUX2_X1 $T=70160 73800 1 0 $X=70045 $Y=72285
X1851 56 46 21 265 52 46 NAND2_X1 $T=20570 68200 0 0 $X=20455 $Y=68085
X1852 57 46 106 107 52 46 NAND2_X1 $T=21900 73800 0 180 $X=21215 $Y=72285
X1853 88 46 86 266 52 46 NAND2_X1 $T=24750 71000 1 180 $X=24065 $Y=70885
X1854 89 46 203 202 52 46 NAND2_X1 $T=25510 71000 1 0 $X=25395 $Y=69485
X1855 91 46 62 254 52 46 NAND2_X1 $T=31970 71000 0 0 $X=31855 $Y=70885
X1856 64 46 112 25 52 46 NAND2_X1 $T=36340 73800 1 0 $X=36225 $Y=72285
X1857 113 46 67 26 52 46 NAND2_X1 $T=40330 73800 1 0 $X=40215 $Y=72285
X1858 261 52 79 104 46 46 NOR2_X1 $T=3090 73800 1 0 $X=2975 $Y=72285
X1859 81 52 82 196 46 46 NOR2_X1 $T=5370 71000 1 180 $X=4685 $Y=70885
X1860 241 52 242 224 46 46 NOR2_X1 $T=13920 71000 0 0 $X=13805 $Y=70885
X1861 245 52 243 244 46 46 NOR2_X1 $T=17150 68200 1 180 $X=16465 $Y=68085
X1862 224 52 244 147 46 46 NOR2_X1 $T=16960 71000 0 0 $X=16845 $Y=70885
X1863 53 52 147 199 46 46 NOR2_X1 $T=18290 73800 0 180 $X=17605 $Y=72285
X1864 19 52 20 246 46 46 NOR2_X1 $T=18670 71000 0 0 $X=18555 $Y=70885
X1865 106 52 246 247 46 46 NOR2_X1 $T=20000 71000 1 0 $X=19885 $Y=69485
X1866 229 52 246 84 46 46 NOR2_X1 $T=20570 71000 1 180 $X=19885 $Y=70885
X1867 55 52 108 83 46 46 NOR2_X1 $T=20190 73800 1 0 $X=20075 $Y=72285
X1868 157 52 55 85 46 46 NOR2_X1 $T=21330 73800 0 180 $X=20645 $Y=72285
X1869 88 52 86 108 46 46 NOR2_X1 $T=22850 73800 0 180 $X=22165 $Y=72285
X1870 89 52 203 267 46 46 NOR2_X1 $T=26080 71000 0 0 $X=25965 $Y=70885
X1871 206 52 251 252 46 46 NOR2_X1 $T=29310 71000 0 0 $X=29195 $Y=70885
X1872 254 52 252 253 46 46 NOR2_X1 $T=31400 71000 1 180 $X=30715 $Y=70885
X1873 269 52 252 148 46 46 NOR2_X1 $T=30830 73800 1 0 $X=30715 $Y=72285
X1874 91 52 62 207 46 46 NOR2_X1 $T=33300 71000 0 0 $X=33185 $Y=70885
X1875 63 52 207 149 46 46 NOR2_X1 $T=34250 73800 1 0 $X=34135 $Y=72285
X1876 64 52 112 24 46 46 NOR2_X1 $T=36340 73800 0 180 $X=35655 $Y=72285
X1877 113 52 67 93 46 46 NOR2_X1 $T=40330 73800 0 180 $X=39645 $Y=72285
X1878 237 52 39 220 46 46 NOR2_X1 $T=70730 68200 0 0 $X=70615 $Y=68085
X1879 101 52 258 221 46 46 NOR2_X1 $T=72060 68200 0 0 $X=71945 $Y=68085
X1880 74 52 258 240 46 46 NOR2_X1 $T=74150 71000 0 180 $X=73465 $Y=69485
X1881 260 52 74 282 46 46 NOR2_X1 $T=75480 71000 1 0 $X=75365 $Y=69485
X1882 42 52 76 258 46 46 NOR2_X1 $T=76810 68200 1 180 $X=76125 $Y=68085
X1883 56 21 200 22 46 52 46 AOI21_X1 $T=21900 68200 1 180 $X=21025 $Y=68085
X1884 266 202 249 231 46 52 46 AOI21_X1 $T=24750 71000 0 0 $X=24635 $Y=70885
X1885 202 204 110 267 46 52 46 AOI21_X1 $T=27600 73800 0 180 $X=26725 $Y=72285
X1886 25 26 268 270 46 52 46 AOI21_X1 $T=36910 73800 1 0 $X=36795 $Y=72285
X1887 237 39 155 290 46 52 46 AOI21_X1 $T=69970 68200 0 0 $X=69855 $Y=68085
X1888 237 39 281 220 46 52 46 AOI21_X1 $T=70350 71000 1 0 $X=70235 $Y=69485
X1889 204 52 267 231 46 250 46 NOR3_X1 $T=26840 73800 0 180 $X=25965 $Y=72285
X1890 66 52 93 270 46 272 46 NOR3_X1 $T=39000 73800 1 0 $X=38885 $Y=72285
X1891 258 52 74 220 46 119 46 NOR3_X1 $T=74150 68200 1 180 $X=73275 $Y=68085
X1892 46 284 261 196 52 46 XNOR2_X1 $T=2330 71000 0 0 $X=2215 $Y=70885
X1893 46 82 262 81 52 46 XNOR2_X1 $T=6510 71000 1 180 $X=5255 $Y=70885
X1894 46 248 58 200 52 46 XNOR2_X1 $T=23420 71000 0 180 $X=22165 $Y=69485
X1895 46 60 59 201 52 46 XNOR2_X1 $T=23610 68200 0 0 $X=23495 $Y=68085
X1896 46 281 156 291 52 46 XNOR2_X1 $T=69970 71000 0 0 $X=69855 $Y=70885
X1897 46 282 169 239 52 46 XNOR2_X1 $T=75290 71000 0 0 $X=75175 $Y=70885
X1898 252 207 24 46 52 270 OR3_X1 $T=34820 73800 1 0 $X=34705 $Y=72285
X1899 110 87 46 109 86 88 52 OAI22_X1 $T=24750 73800 0 180 $X=23685 $Y=72285
X1900 259 101 46 239 76 42 52 OAI22_X1 $T=75290 68200 0 0 $X=75175 $Y=68085
X1901 250 52 249 247 229 248 46 46 NOR4_X1 $T=23040 71000 1 180 $X=21975 $Y=70885
X1902 272 52 268 253 269 204 46 46 NOR4_X1 $T=29880 73800 1 0 $X=29765 $Y=72285
X1903 284 4 262 263 52 46 47 46 FA_X1 $T=3660 73800 1 0 $X=3545 $Y=72285
X1904 203 173 90 174 52 46 206 46 FA_X1 $T=25700 68200 0 0 $X=25585 $Y=68085
X1905 251 205 111 158 52 46 91 46 FA_X1 $T=26840 71000 1 0 $X=26725 $Y=69485
X1906 205 23 92 159 52 46 208 46 FA_X1 $T=31590 68200 0 0 $X=31475 $Y=68085
X1907 62 208 271 122 52 46 64 46 FA_X1 $T=35770 71000 1 0 $X=35655 $Y=69485
X1908 112 209 255 65 52 46 113 46 FA_X1 $T=35770 71000 0 0 $X=35655 $Y=70885
X1909 271 232 163 160 52 46 209 46 FA_X1 $T=38810 71000 1 0 $X=38695 $Y=69485
X1910 255 210 94 175 52 46 133 46 FA_X1 $T=38810 71000 0 0 $X=38695 $Y=70885
X1911 232 27 95 123 52 46 134 46 FA_X1 $T=40140 68200 0 0 $X=40025 $Y=68085
X1912 150 211 124 125 52 46 212 46 FA_X1 $T=45270 71000 1 180 $X=42115 $Y=70885
X1913 210 170 126 140 52 46 286 46 FA_X1 $T=43180 68200 0 0 $X=43065 $Y=68085
X1914 211 127 114 274 52 46 273 46 FA_X1 $T=46410 71000 1 0 $X=46295 $Y=69485
X1915 151 212 233 286 52 46 135 46 FA_X1 $T=46980 73800 1 0 $X=46865 $Y=72285
X1916 233 287 171 128 52 46 215 46 FA_X1 $T=49830 71000 0 0 $X=49715 $Y=70885
X1917 274 172 256 164 52 46 214 46 FA_X1 $T=50210 68200 0 0 $X=50095 $Y=68085
X1918 287 214 72 276 52 46 275 46 FA_X1 $T=52870 71000 0 0 $X=52755 $Y=70885
X1919 152 215 273 294 52 46 136 46 FA_X1 $T=53440 73800 1 0 $X=53325 $Y=72285
X1920 256 31 97 161 52 46 236 46 FA_X1 $T=55910 68200 0 0 $X=55795 $Y=68085
X1921 153 216 277 275 52 46 115 46 FA_X1 $T=57620 73800 1 0 $X=57505 $Y=72285
X1922 217 32 98 165 52 46 278 46 FA_X1 $T=58950 68200 0 0 $X=58835 $Y=68085
X1923 294 217 176 288 52 46 216 46 FA_X1 $T=58950 71000 1 0 $X=58835 $Y=69485
X1924 276 166 99 236 52 46 289 46 FA_X1 $T=59710 71000 0 0 $X=59595 $Y=70885
X1925 288 177 178 162 52 46 257 46 FA_X1 $T=62370 71000 1 0 $X=62255 $Y=69485
X1926 277 283 257 289 52 46 218 46 FA_X1 $T=62750 71000 0 0 $X=62635 $Y=70885
X1927 116 218 117 278 52 46 237 46 FA_X1 $T=65410 71000 1 0 $X=65295 $Y=69485
X1928 283 38 100 168 52 46 139 46 FA_X1 $T=69970 68200 1 180 $X=66815 $Y=68085
X1930 118 46 221 41 52 238 NAND3_X1 $T=72820 71000 1 0 $X=72705 $Y=69485
X1932 198 46 52 105 CLKBUF_X1 $T=15250 71000 0 180 $X=14565 $Y=69485
X1933 264 46 52 54 CLKBUF_X1 $T=18670 71000 1 0 $X=18555 $Y=69485
X1934 224 51 52 199 18 46 244 264 AOI221_X1 $T=17530 71000 0 0 $X=17415 $Y=70885
X1935 81 5 6 8 46 52 228 OR4_X1 $T=9550 71000 1 0 $X=9435 $Y=69485
X1936 197 7 9 10 46 52 223 OR4_X1 $T=10690 71000 1 0 $X=10575 $Y=69485
X1937 82 12 13 14 46 52 226 OR4_X1 $T=13540 71000 1 0 $X=13425 $Y=69485
X1938 50 15 16 17 46 52 227 OR4_X1 $T=15820 71000 1 0 $X=15705 $Y=69485
X1939 8 46 6 5 81 245 52 NAND4_X1 $T=8410 68200 0 0 $X=8295 $Y=68085
X1940 9 46 7 197 82 241 52 NAND4_X1 $T=10690 71000 0 0 $X=10575 $Y=70885
X1941 14 46 13 12 10 242 52 NAND4_X1 $T=13920 71000 1 180 $X=12855 $Y=70885
X1942 17 46 16 15 50 243 52 NAND4_X1 $T=16580 68200 1 180 $X=15515 $Y=68085
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
** N=279 EP=180 IP=2365 FDC=1514
X1173 138 2 24 23 142 DFF_X1 $T=1000 65400 1 0 $X=885 $Y=63885
X1174 139 2 24 23 25 DFF_X1 $T=2330 65400 0 0 $X=2215 $Y=65285
X1175 267 2 24 23 26 DFF_X1 $T=4800 68200 1 0 $X=4685 $Y=66685
X1176 28 2 24 23 143 DFF_X1 $T=12020 65400 1 0 $X=11905 $Y=63885
X1177 268 2 24 23 144 DFF_X1 $T=12400 68200 1 0 $X=12285 $Y=66685
X1178 140 8 24 23 110 DFF_X1 $T=15630 65400 0 0 $X=15515 $Y=65285
X1179 145 8 24 23 146 DFF_X1 $T=18860 68200 0 180 $X=15515 $Y=66685
X1180 228 2 24 23 77 DFF_X1 $T=18670 65400 1 0 $X=18555 $Y=63885
X1181 19 20 24 23 137 DFF_X1 $T=78710 68200 1 0 $X=78595 $Y=66685
X1182 22 1 24 23 108 24 AND2_X1 $T=1190 68200 1 0 $X=1075 $Y=66685
X1183 22 3 24 23 73 24 AND2_X1 $T=2330 68200 1 0 $X=2215 $Y=66685
X1184 22 4 24 23 267 24 AND2_X1 $T=4040 68200 1 0 $X=3925 $Y=66685
X1185 22 5 24 23 109 24 AND2_X1 $T=8030 62600 0 0 $X=7915 $Y=62485
X1186 22 6 24 23 268 24 AND2_X1 $T=10500 65400 0 180 $X=9625 $Y=63885
X1187 22 7 24 23 228 24 AND2_X1 $T=11450 65400 0 0 $X=11335 $Y=65285
X1314 51 18 255 256 24 23 OAI21_X1 $T=70730 65400 0 0 $X=70615 $Y=65285
X1315 51 18 86 52 24 23 OAI21_X1 $T=71490 65400 1 0 $X=71375 $Y=63885
X1316 156 243 128 52 24 23 OAI21_X1 $T=72630 68200 1 0 $X=72515 $Y=66685
X1363 256 24 23 243 24 INV_X1 $T=72630 65400 0 180 $X=72135 $Y=63885
X1488 35 40 24 23 INV_X2 $T=36340 62600 0 0 $X=36225 $Y=62485
X1489 44 63 24 23 INV_X2 $T=43370 62600 0 0 $X=43255 $Y=62485
X1490 14 15 24 23 INV_X2 $T=45270 65400 0 0 $X=45155 $Y=65285
X1491 62 64 24 23 INV_X2 $T=46980 65400 1 0 $X=46865 $Y=63885
X1492 13 46 24 23 INV_X2 $T=48880 65400 1 0 $X=48765 $Y=63885
X1493 61 81 24 23 INV_X2 $T=51920 65400 1 0 $X=51805 $Y=63885
X1494 66 68 24 23 INV_X2 $T=57240 62600 0 0 $X=57125 $Y=62485
X1540 74 24 257 147 23 24 NAND2_X1 $T=18860 68200 1 0 $X=18745 $Y=66685
X1541 51 24 18 256 23 24 NAND2_X1 $T=70920 65400 1 0 $X=70805 $Y=63885
X1542 242 24 265 89 23 24 NAND2_X1 $T=75860 68200 1 0 $X=75745 $Y=66685
X1543 74 23 257 148 24 24 NOR2_X1 $T=19430 68200 1 0 $X=19315 $Y=66685
X1544 75 23 76 30 24 24 NOR2_X1 $T=20760 68200 1 0 $X=20645 $Y=66685
X1545 57 23 33 58 24 24 NOR2_X1 $T=35010 62600 0 0 $X=34895 $Y=62485
X1546 57 23 41 246 24 24 NOR2_X1 $T=38430 62600 0 0 $X=38315 $Y=62485
X1547 40 23 33 247 24 24 NOR2_X1 $T=39570 62600 1 180 $X=38885 $Y=62485
X1548 40 23 41 248 24 24 NOR2_X1 $T=41280 62600 0 0 $X=41165 $Y=62485
X1549 15 23 33 240 24 24 NOR2_X1 $T=43370 62600 1 180 $X=42685 $Y=62485
X1550 15 23 41 241 24 24 NOR2_X1 $T=45460 65400 1 0 $X=45345 $Y=63885
X1551 63 23 33 261 24 24 NOR2_X1 $T=48120 62600 1 180 $X=47435 $Y=62485
X1552 63 23 41 232 24 24 NOR2_X1 $T=49070 62600 0 0 $X=48955 $Y=62485
X1553 64 23 33 263 24 24 NOR2_X1 $T=50210 65400 1 0 $X=50095 $Y=63885
X1554 64 23 41 234 24 24 NOR2_X1 $T=54010 62600 0 0 $X=53895 $Y=62485
X1555 46 23 33 250 24 24 NOR2_X1 $T=55530 62600 0 0 $X=55415 $Y=62485
X1556 40 23 161 133 24 24 NOR2_X1 $T=56100 62600 0 0 $X=55985 $Y=62485
X1557 15 23 70 65 24 24 NOR2_X1 $T=56670 62600 0 0 $X=56555 $Y=62485
X1558 46 23 41 236 24 24 NOR2_X1 $T=58760 62600 0 0 $X=58645 $Y=62485
X1559 81 23 33 251 24 24 NOR2_X1 $T=59900 65400 1 0 $X=59785 $Y=63885
X1560 63 23 70 134 24 24 NOR2_X1 $T=60090 62600 0 0 $X=59975 $Y=62485
X1561 64 23 71 135 24 24 NOR2_X1 $T=61420 62600 0 0 $X=61305 $Y=62485
X1562 68 23 33 136 24 24 NOR2_X1 $T=65030 62600 0 0 $X=64915 $Y=62485
X1563 63 23 161 238 24 24 NOR2_X1 $T=67120 62600 0 0 $X=67005 $Y=62485
X1564 64 23 70 253 24 24 NOR2_X1 $T=68260 62600 1 180 $X=67575 $Y=62485
X1565 46 23 71 254 24 24 NOR2_X1 $T=68830 62600 1 180 $X=68145 $Y=62485
X1566 242 23 265 129 24 24 NOR2_X1 $T=77000 68200 0 180 $X=76315 $Y=66685
X1567 24 87 50 255 23 24 XNOR2_X1 $T=68450 65400 0 0 $X=68335 $Y=65285
X1568 87 243 24 180 18 51 23 OAI22_X1 $T=72630 68200 0 180 $X=71565 $Y=66685
X1569 42 23 13 44 14 102 24 24 NOR4_X1 $T=44510 65400 1 0 $X=44395 $Y=63885
X1570 66 23 61 62 35 122 24 24 NOR4_X1 $T=45840 65400 0 0 $X=45725 $Y=65285
X1571 29 91 56 93 23 24 75 24 FA_X1 $T=18860 62600 0 0 $X=18745 $Y=62485
X1572 257 92 244 157 23 24 111 24 FA_X1 $T=18860 65400 0 0 $X=18745 $Y=65285
X1573 244 9 78 167 23 24 269 24 FA_X1 $T=22280 65400 1 0 $X=22165 $Y=63885
X1574 245 229 168 258 23 24 112 24 FA_X1 $T=25320 65400 1 180 $X=22165 $Y=65285
X1575 113 269 245 275 23 24 141 24 FA_X1 $T=22280 68200 1 0 $X=22165 $Y=66685
X1576 275 10 31 169 23 24 114 24 FA_X1 $T=25320 65400 1 0 $X=25205 $Y=63885
X1577 258 277 182 95 23 24 270 24 FA_X1 $T=28360 65400 1 0 $X=28245 $Y=63885
X1578 149 276 32 270 23 24 115 24 FA_X1 $T=28740 68200 1 0 $X=28625 $Y=66685
X1579 229 11 170 94 23 24 116 24 FA_X1 $T=28930 62600 0 0 $X=28815 $Y=62485
X1580 276 271 259 171 23 24 117 24 FA_X1 $T=31400 65400 1 0 $X=31285 $Y=63885
X1581 277 96 97 158 23 24 271 24 FA_X1 $T=31970 62600 0 0 $X=31855 $Y=62485
X1582 259 98 172 272 23 24 230 24 FA_X1 $T=33490 65400 0 0 $X=33375 $Y=65285
X1583 150 12 34 99 23 24 118 24 FA_X1 $T=37480 65400 0 180 $X=34325 $Y=63885
X1584 151 230 21 37 23 24 119 24 FA_X1 $T=38810 68200 0 180 $X=35655 $Y=66685
X1585 272 246 247 14 23 24 266 24 FA_X1 $T=37480 65400 1 0 $X=37365 $Y=63885
X1586 152 38 266 159 23 24 59 24 FA_X1 $T=41850 68200 0 180 $X=38695 $Y=66685
X1587 36 248 240 44 23 24 231 24 FA_X1 $T=40520 65400 1 0 $X=40405 $Y=63885
X1588 120 231 43 101 23 24 60 24 FA_X1 $T=42230 65400 0 0 $X=42115 $Y=65285
X1589 79 100 260 39 23 24 121 24 FA_X1 $T=45270 68200 0 180 $X=42115 $Y=66685
X1590 131 241 261 62 23 24 260 24 FA_X1 $T=43940 62600 0 0 $X=43825 $Y=62485
X1591 132 232 263 13 23 24 45 24 FA_X1 $T=46790 65400 0 0 $X=46675 $Y=65285
X1592 80 262 173 160 23 24 55 24 FA_X1 $T=49070 68200 1 0 $X=48955 $Y=66685
X1593 262 16 176 249 23 24 233 24 FA_X1 $T=49640 62600 0 0 $X=49525 $Y=62485
X1594 153 233 53 278 23 24 47 24 FA_X1 $T=52110 68200 1 0 $X=51995 $Y=66685
X1595 249 234 250 61 23 24 235 24 FA_X1 $T=55910 65400 0 0 $X=55795 $Y=65285
X1596 278 235 82 162 23 24 123 24 FA_X1 $T=56860 65400 1 0 $X=56745 $Y=63885
X1597 67 236 251 66 23 24 273 24 FA_X1 $T=58950 65400 0 0 $X=58835 $Y=65285
X1598 48 49 103 174 23 24 124 24 FA_X1 $T=62370 65400 1 0 $X=62255 $Y=63885
X1599 83 17 252 179 23 24 237 24 FA_X1 $T=62370 65400 0 0 $X=62255 $Y=65285
X1600 154 237 84 273 23 24 125 24 FA_X1 $T=63510 68200 1 0 $X=63395 $Y=66685
X1601 252 238 253 254 23 24 126 24 FA_X1 $T=65410 65400 1 0 $X=65295 $Y=63885
X1602 69 105 104 163 23 24 127 24 FA_X1 $T=65410 65400 0 0 $X=65295 $Y=65285
X1603 155 106 72 177 23 24 264 24 FA_X1 $T=68830 62600 0 0 $X=68715 $Y=62485
X1604 85 274 279 164 23 24 242 24 FA_X1 $T=71490 65400 0 0 $X=71375 $Y=65285
X1605 88 181 264 175 23 24 274 24 FA_X1 $T=75670 65400 0 180 $X=72515 $Y=63885
X1606 279 178 107 165 23 24 239 24 FA_X1 $T=78900 62600 0 0 $X=78785 $Y=62485
X1607 265 239 90 166 23 24 130 24 FA_X1 $T=81370 65400 1 0 $X=81255 $Y=63885
.ENDS
***************************************
.SUBCKT ICV_14
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=2 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 VSS VDD ZN
** N=11 EP=7 IP=0 FDC=10
M0 9 A1 8 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 10 A2 9 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 11 A3 10 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 11 VSS NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 8 VSS VSS NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 8 A1 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD A2 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 8 A3 VDD VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 8 VDD PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 8 VDD VDD PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 94 95 97 98 99 100 101 102 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163 164
+ 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183 184
+ 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203 204
+ 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219
** N=419 EP=215 IP=5466 FDC=3022
X2633 26 7 33 26 130 DFF_X1 $T=2330 57000 1 0 $X=2215 $Y=55485
X2634 349 7 33 26 101 DFF_X1 $T=2330 57000 0 0 $X=2215 $Y=56885
X2635 303 7 33 26 41 DFF_X1 $T=3090 59800 1 0 $X=2975 $Y=58285
X2636 348 7 33 26 169 DFF_X1 $T=4420 54200 0 0 $X=4305 $Y=54085
X2637 245 12 33 26 102 DFF_X1 $T=5180 62600 1 0 $X=5065 $Y=61085
X2638 246 7 33 26 249 DFF_X1 $T=7650 54200 0 0 $X=7535 $Y=54085
X2639 396 7 33 26 43 DFF_X1 $T=7650 57000 1 0 $X=7535 $Y=55485
X2640 304 12 33 26 131 DFF_X1 $T=8030 51400 0 0 $X=7915 $Y=51285
X2641 397 7 33 26 103 DFF_X1 $T=12590 59800 0 0 $X=12475 $Y=59685
X2642 306 12 33 26 301 DFF_X1 $T=13540 59800 1 0 $X=13425 $Y=58285
X2643 305 7 33 26 277 DFF_X1 $T=13730 54200 1 0 $X=13615 $Y=52685
X2644 100 12 33 26 104 DFF_X1 $T=14300 62600 1 0 $X=14185 $Y=61085
X2645 398 7 33 26 133 DFF_X1 $T=15060 57000 1 0 $X=14945 $Y=55485
X2646 195 7 33 26 144 DFF_X1 $T=53440 51400 0 0 $X=53325 $Y=51285
X2694 38 1 33 26 348 33 AND2_X1 $T=1000 54200 0 0 $X=885 $Y=54085
X2695 38 2 33 26 26 33 AND2_X1 $T=1190 54200 1 0 $X=1075 $Y=52685
X2696 37 3 33 26 245 33 AND2_X1 $T=2710 59800 1 180 $X=1835 $Y=59685
X2697 37 4 33 26 39 33 AND2_X1 $T=2330 51400 0 0 $X=2215 $Y=51285
X2698 38 5 33 26 303 33 AND2_X1 $T=2330 59800 1 0 $X=2215 $Y=58285
X2699 37 6 33 26 40 33 AND2_X1 $T=2330 62600 1 0 $X=2215 $Y=61085
X2700 38 99 33 26 349 33 AND2_X1 $T=3660 54200 0 0 $X=3545 $Y=54085
X2701 38 8 33 26 246 33 AND2_X1 $T=3850 51400 0 0 $X=3735 $Y=51285
X2702 37 9 33 26 167 33 AND2_X1 $T=4420 62600 1 0 $X=4305 $Y=61085
X2703 37 10 33 26 196 33 AND2_X1 $T=5180 59800 0 0 $X=5065 $Y=59685
X2704 37 11 33 26 168 33 AND2_X1 $T=6510 51400 1 180 $X=5635 $Y=51285
X2705 38 13 33 26 396 33 AND2_X1 $T=6700 54200 1 0 $X=6585 $Y=52685
X2706 38 14 33 26 397 33 AND2_X1 $T=6890 57000 1 0 $X=6775 $Y=55485
X2707 37 15 33 26 304 33 AND2_X1 $T=7270 51400 0 0 $X=7155 $Y=51285
X2708 38 16 33 26 197 33 AND2_X1 $T=8600 59800 1 180 $X=7725 $Y=59685
X2709 38 17 33 26 42 33 AND2_X1 $T=8600 59800 0 0 $X=8485 $Y=59685
X2710 38 18 33 26 398 33 AND2_X1 $T=9930 57000 0 0 $X=9815 $Y=56885
X2711 38 19 33 26 305 33 AND2_X1 $T=10120 54200 1 0 $X=10005 $Y=52685
X2712 37 20 33 26 306 33 AND2_X1 $T=10690 59800 1 0 $X=10575 $Y=58285
X3087 133 33 26 85 33 INV_X1 $T=23230 57000 1 0 $X=23115 $Y=55485
X3354 249 90 33 26 INV_X2 $T=14300 54200 0 0 $X=14185 $Y=54085
X3355 22 64 33 26 INV_X2 $T=17530 54200 0 180 $X=16845 $Y=52685
X3356 277 49 33 26 INV_X2 $T=19620 54200 1 0 $X=19505 $Y=52685
X3357 104 50 33 26 INV_X2 $T=19810 59800 1 0 $X=19695 $Y=58285
X3358 135 52 33 26 INV_X2 $T=21140 54200 1 0 $X=21025 $Y=52685
X3359 131 54 33 26 INV_X2 $T=23610 51400 0 0 $X=23495 $Y=51285
X3360 137 30 33 26 INV_X2 $T=24370 57000 1 0 $X=24255 $Y=55485
X3361 106 60 33 26 INV_X2 $T=25510 57000 1 180 $X=24825 $Y=56885
X3362 301 76 33 26 INV_X2 $T=25130 51400 0 0 $X=25015 $Y=51285
X3363 138 63 33 26 INV_X2 $T=29880 59800 1 0 $X=29765 $Y=58285
X3364 140 68 33 26 INV_X2 $T=38240 54200 1 0 $X=38125 $Y=52685
X3365 72 87 33 26 INV_X2 $T=42800 54200 0 0 $X=42685 $Y=54085
X3366 26 124 33 26 INV_X2 $T=43370 54200 0 0 $X=43255 $Y=54085
X3367 81 193 33 26 INV_X2 $T=58380 51400 0 0 $X=58265 $Y=51285
X3461 26 183 200 184 33 33 XOR2_X1 $T=57240 51400 0 0 $X=57125 $Y=51285
X3464 49 26 50 350 33 33 NOR2_X1 $T=19620 54200 0 0 $X=19505 $Y=54085
X3465 85 26 52 247 33 33 NOR2_X1 $T=21900 54200 1 180 $X=21215 $Y=54085
X3466 85 26 50 399 33 33 NOR2_X1 $T=21900 57000 0 180 $X=21215 $Y=55485
X3467 59 26 52 250 33 33 NOR2_X1 $T=21330 59800 1 0 $X=21215 $Y=58285
X3468 85 26 54 353 33 33 NOR2_X1 $T=23610 51400 1 180 $X=22925 $Y=51285
X3469 55 26 50 309 33 33 NOR2_X1 $T=23800 57000 1 180 $X=23115 $Y=56885
X3470 85 26 24 354 33 33 NOR2_X1 $T=23800 57000 1 0 $X=23685 $Y=55485
X3471 64 26 54 310 33 33 NOR2_X1 $T=24940 57000 1 0 $X=24825 $Y=55485
X3472 49 26 76 251 33 33 NOR2_X1 $T=26270 54200 0 180 $X=25585 $Y=52685
X3473 55 26 52 253 33 33 NOR2_X1 $T=26270 59800 1 0 $X=26155 $Y=58285
X3474 49 26 24 279 33 33 NOR2_X1 $T=27030 54200 0 0 $X=26915 $Y=54085
X3475 90 26 50 378 33 33 NOR2_X1 $T=28550 59800 0 180 $X=27865 $Y=58285
X3476 59 26 54 313 33 33 NOR2_X1 $T=28740 54200 1 180 $X=28055 $Y=54085
X3477 85 26 63 280 33 33 NOR2_X1 $T=29310 54200 0 180 $X=28625 $Y=52685
X3478 64 26 76 355 33 33 NOR2_X1 $T=29880 57000 0 180 $X=29195 $Y=55485
X3479 85 26 60 356 33 33 NOR2_X1 $T=29880 57000 1 180 $X=29195 $Y=56885
X3480 49 26 60 357 33 33 NOR2_X1 $T=30070 51400 1 180 $X=29385 $Y=51285
X3481 90 26 52 281 33 33 NOR2_X1 $T=31590 57000 1 180 $X=30905 $Y=56885
X3482 64 26 24 315 33 33 NOR2_X1 $T=31210 51400 0 0 $X=31095 $Y=51285
X3483 85 26 65 254 33 33 NOR2_X1 $T=31590 57000 0 0 $X=31475 $Y=56885
X3484 30 26 50 314 33 33 NOR2_X1 $T=32350 59800 0 180 $X=31665 $Y=58285
X3485 59 26 76 358 33 33 NOR2_X1 $T=32920 54200 0 180 $X=32235 $Y=52685
X3486 30 26 52 255 33 33 NOR2_X1 $T=33490 59800 1 0 $X=33375 $Y=58285
X3487 49 26 63 360 33 33 NOR2_X1 $T=34630 54200 0 0 $X=34515 $Y=54085
X3488 85 26 68 316 33 33 NOR2_X1 $T=35010 54200 1 0 $X=34895 $Y=52685
X3489 59 26 24 401 33 33 NOR2_X1 $T=35010 59800 1 0 $X=34895 $Y=58285
X3490 64 26 60 380 33 33 NOR2_X1 $T=35580 57000 1 0 $X=35465 $Y=55485
X3491 55 26 76 402 33 33 NOR2_X1 $T=37100 57000 1 180 $X=36415 $Y=56885
X3492 90 26 54 414 33 33 NOR2_X1 $T=37290 59800 0 180 $X=36605 $Y=58285
X3493 49 26 65 256 33 33 NOR2_X1 $T=38240 51400 0 0 $X=38125 $Y=51285
X3494 55 26 24 257 33 33 NOR2_X1 $T=38240 57000 0 0 $X=38125 $Y=56885
X3495 90 26 24 403 33 33 NOR2_X1 $T=38430 59800 1 0 $X=38315 $Y=58285
X3496 90 26 76 361 33 33 NOR2_X1 $T=39570 57000 1 0 $X=39455 $Y=55485
X3497 30 26 76 362 33 33 NOR2_X1 $T=40520 59800 0 180 $X=39835 $Y=58285
X3498 30 26 54 363 33 33 NOR2_X1 $T=40140 57000 1 0 $X=40025 $Y=55485
X3499 86 26 54 364 33 33 NOR2_X1 $T=40330 62600 1 0 $X=40215 $Y=61085
X3500 64 26 65 319 33 33 NOR2_X1 $T=42800 57000 0 0 $X=42685 $Y=56885
X3501 59 26 63 320 33 33 NOR2_X1 $T=43370 57000 0 0 $X=43255 $Y=56885
X3502 55 26 60 321 33 33 NOR2_X1 $T=45460 57000 1 180 $X=44775 $Y=56885
X3503 30 26 24 323 33 33 NOR2_X1 $T=45270 54200 1 0 $X=45155 $Y=52685
X3504 86 26 76 324 33 33 NOR2_X1 $T=48120 54200 0 180 $X=47435 $Y=52685
X3505 95 26 54 260 33 33 NOR2_X1 $T=48310 54200 1 180 $X=47625 $Y=54085
X3506 55 26 65 386 33 33 NOR2_X1 $T=48880 57000 0 180 $X=48195 $Y=55485
X3507 90 26 63 325 33 33 NOR2_X1 $T=49640 54200 1 180 $X=48955 $Y=54085
X3508 86 26 24 302 33 33 NOR2_X1 $T=49260 59800 1 0 $X=49145 $Y=58285
X3509 30 26 60 326 33 33 NOR2_X1 $T=50210 54200 1 180 $X=49525 $Y=54085
X3510 95 26 76 385 33 33 NOR2_X1 $T=50400 59800 1 0 $X=50285 $Y=58285
X3511 85 26 75 286 33 33 NOR2_X1 $T=51350 51400 1 180 $X=50665 $Y=51285
X3512 79 26 54 417 33 33 NOR2_X1 $T=50970 59800 1 0 $X=50855 $Y=58285
X3513 49 26 87 327 33 33 NOR2_X1 $T=51920 54200 0 0 $X=51805 $Y=54085
X3514 49 26 78 261 33 33 NOR2_X1 $T=51920 57000 1 0 $X=51805 $Y=55485
X3515 64 26 83 288 33 33 NOR2_X1 $T=54010 54200 1 180 $X=53325 $Y=54085
X3516 59 26 68 328 33 33 NOR2_X1 $T=53630 57000 1 0 $X=53515 $Y=55485
X3517 64 26 78 262 33 33 NOR2_X1 $T=54010 54200 0 0 $X=53895 $Y=54085
X3518 90 26 65 388 33 33 NOR2_X1 $T=55340 57000 1 0 $X=55225 $Y=55485
X3519 59 26 83 331 33 33 NOR2_X1 $T=57240 51400 1 180 $X=56555 $Y=51285
X3520 86 26 60 367 33 33 NOR2_X1 $T=56670 59800 1 0 $X=56555 $Y=58285
X3521 126 26 54 290 33 33 NOR2_X1 $T=57050 62600 1 0 $X=56935 $Y=61085
X3522 55 26 68 405 33 33 NOR2_X1 $T=58000 54200 0 180 $X=57315 $Y=52685
X3523 30 26 63 330 33 33 NOR2_X1 $T=58000 57000 1 180 $X=57315 $Y=56885
X3524 79 26 24 332 33 33 NOR2_X1 $T=59330 59800 0 0 $X=59215 $Y=59685
X3525 59 26 78 368 33 33 NOR2_X1 $T=59710 57000 1 0 $X=59595 $Y=55485
X3526 55 26 83 292 33 33 NOR2_X1 $T=60280 54200 0 0 $X=60165 $Y=54085
X3527 90 26 68 333 33 33 NOR2_X1 $T=61420 57000 1 0 $X=61305 $Y=55485
X3528 30 26 65 266 33 33 NOR2_X1 $T=62180 57000 0 0 $X=62065 $Y=56885
X3529 146 26 52 267 33 33 NOR2_X1 $T=62370 62600 1 0 $X=62255 $Y=61085
X3530 49 26 124 335 33 33 NOR2_X1 $T=63130 51400 0 0 $X=63015 $Y=51285
X3531 86 26 63 337 33 33 NOR2_X1 $T=64080 59800 0 180 $X=63395 $Y=58285
X3532 85 26 124 265 33 33 NOR2_X1 $T=63700 54200 0 0 $X=63585 $Y=54085
X3533 95 26 60 336 33 33 NOR2_X1 $T=63700 57000 0 0 $X=63585 $Y=56885
X3534 59 26 87 338 33 33 NOR2_X1 $T=65220 51400 1 180 $X=64535 $Y=51285
X3535 64 26 75 370 33 33 NOR2_X1 $T=65410 54200 0 180 $X=64725 $Y=52685
X3536 49 26 75 294 33 33 NOR2_X1 $T=66550 54200 0 180 $X=65865 $Y=52685
X3537 64 26 87 339 33 33 NOR2_X1 $T=65980 54200 0 0 $X=65865 $Y=54085
X3538 86 26 65 268 33 33 NOR2_X1 $T=65980 59800 1 0 $X=65865 $Y=58285
X3539 55 26 78 341 33 33 NOR2_X1 $T=67690 54200 1 0 $X=67575 $Y=52685
X3540 95 26 65 269 33 33 NOR2_X1 $T=68260 57000 0 180 $X=67575 $Y=55485
X3541 95 26 63 371 33 33 NOR2_X1 $T=68070 59800 1 0 $X=67955 $Y=58285
X3542 79 26 60 391 33 33 NOR2_X1 $T=68640 59800 1 0 $X=68525 $Y=58285
X3543 90 26 83 407 33 33 NOR2_X1 $T=69780 54200 0 180 $X=69095 $Y=52685
X3544 126 26 60 419 33 33 NOR2_X1 $T=70540 57000 1 180 $X=69855 $Y=56885
X3545 79 26 63 411 33 33 NOR2_X1 $T=71110 57000 1 180 $X=70425 $Y=56885
X3546 30 26 68 296 33 33 NOR2_X1 $T=71300 54200 0 180 $X=70615 $Y=52685
X3547 86 26 68 408 33 33 NOR2_X1 $T=72630 57000 1 0 $X=72515 $Y=55485
X3548 90 26 78 271 33 33 NOR2_X1 $T=73770 57000 0 180 $X=73085 $Y=55485
X3549 30 26 83 298 33 33 NOR2_X1 $T=74530 54200 0 0 $X=74415 $Y=54085
X3550 64 26 124 412 33 33 NOR2_X1 $T=76240 54200 0 0 $X=76125 $Y=54085
X3551 55 26 87 375 33 33 NOR2_X1 $T=78140 54200 0 0 $X=78025 $Y=54085
X3552 59 26 75 376 33 33 NOR2_X1 $T=78330 51400 0 0 $X=78215 $Y=51285
X3554 44 26 48 22 277 318 33 33 NOR4_X1 $T=18670 54200 1 0 $X=18555 $Y=52685
X3555 137 26 249 53 133 352 33 33 NOR4_X1 $T=23230 57000 0 180 $X=22165 $Y=55485
X3556 138 26 106 301 104 57 33 33 NOR4_X1 $T=26270 59800 0 180 $X=25205 $Y=58285
X3557 208 26 26 72 140 191 33 33 NOR4_X1 $T=37290 54200 1 0 $X=37175 $Y=52685
X3558 132 45 307 276 26 33 134 33 FA_X1 $T=15820 59800 0 0 $X=15705 $Y=59685
X3559 276 247 350 22 26 33 278 33 FA_X1 $T=16580 54200 0 0 $X=16465 $Y=54085
X3560 170 21 51 278 26 33 105 33 FA_X1 $T=16770 59800 1 0 $X=16655 $Y=58285
X3561 171 135 399 277 26 33 307 33 FA_X1 $T=18290 57000 1 0 $X=18175 $Y=55485
X3562 46 152 301 353 26 33 136 33 FA_X1 $T=18860 51400 0 0 $X=18745 $Y=51285
X3563 47 248 351 308 26 33 172 33 FA_X1 $T=18860 59800 0 0 $X=18745 $Y=59685
X3564 308 354 251 310 26 33 56 33 FA_X1 $T=21710 54200 1 0 $X=21595 $Y=52685
X3565 351 250 309 249 26 33 23 33 FA_X1 $T=22280 59800 1 0 $X=22165 $Y=58285
X3566 248 252 311 106 26 33 107 33 FA_X1 $T=22850 62600 1 0 $X=22735 $Y=61085
X3567 311 279 355 313 26 33 108 33 FA_X1 $T=25510 57000 1 0 $X=25395 $Y=55485
X3568 58 312 138 356 26 33 173 33 FA_X1 $T=28550 57000 1 180 $X=25395 $Y=56885
X3569 252 253 378 137 26 33 109 33 FA_X1 $T=25510 59800 0 0 $X=25395 $Y=59685
X3570 312 153 280 357 26 33 400 33 FA_X1 $T=25700 51400 0 0 $X=25585 $Y=51285
X3571 198 281 314 44 26 33 174 33 FA_X1 $T=28550 59800 0 0 $X=28435 $Y=59685
X3572 61 315 358 206 26 33 379 33 FA_X1 $T=29310 54200 1 0 $X=29195 $Y=52685
X3573 67 379 400 317 26 33 62 33 FA_X1 $T=32920 57000 0 180 $X=29765 $Y=55485
X3574 69 25 110 316 26 33 359 33 FA_X1 $T=34820 51400 1 180 $X=31665 $Y=51285
X3575 111 254 360 380 26 33 112 33 FA_X1 $T=33490 57000 0 0 $X=33375 $Y=56885
X3576 66 255 139 207 26 33 113 33 FA_X1 $T=34250 62600 1 0 $X=34135 $Y=61085
X3577 141 401 402 414 26 33 175 33 FA_X1 $T=39570 59800 1 180 $X=36415 $Y=59685
X3578 114 154 282 416 26 33 115 33 FA_X1 $T=37290 62600 1 0 $X=37175 $Y=61085
X3579 317 409 381 140 26 33 70 33 FA_X1 $T=40900 54200 1 180 $X=37745 $Y=54085
X3580 381 256 213 217 26 33 365 33 FA_X1 $T=38810 51400 0 0 $X=38695 $Y=51285
X3581 36 365 359 382 26 33 71 33 FA_X1 $T=38810 54200 1 0 $X=38695 $Y=52685
X3582 409 257 361 363 26 33 178 33 FA_X1 $T=38810 57000 0 0 $X=38695 $Y=56885
X3583 282 403 362 364 26 33 179 33 FA_X1 $T=39570 59800 0 0 $X=39455 $Y=59685
X3584 382 384 116 209 26 33 283 33 FA_X1 $T=42230 51400 0 0 $X=42115 $Y=51285
X3585 35 215 283 383 26 33 117 33 FA_X1 $T=42230 57000 1 0 $X=42115 $Y=55485
X3586 416 319 320 321 26 33 118 33 FA_X1 $T=42230 59800 1 0 $X=42115 $Y=58285
X3587 199 27 322 155 26 33 119 33 FA_X1 $T=42230 62600 1 0 $X=42115 $Y=61085
X3588 383 258 218 410 26 33 181 33 FA_X1 $T=43370 59800 0 0 $X=43255 $Y=59685
X3589 384 323 324 260 26 33 143 33 FA_X1 $T=43940 54200 0 0 $X=43825 $Y=54085
X3590 259 386 325 326 26 33 289 33 FA_X1 $T=45270 57000 1 0 $X=45155 $Y=55485
X3591 322 259 284 72 26 33 73 33 FA_X1 $T=45270 59800 1 0 $X=45155 $Y=58285
X3592 410 302 385 417 26 33 285 33 FA_X1 $T=45270 62600 1 0 $X=45155 $Y=61085
X3593 192 26 286 327 26 33 287 33 FA_X1 $T=48120 54200 1 0 $X=48005 $Y=52685
X3594 284 261 288 328 26 33 329 33 FA_X1 $T=51350 57000 0 0 $X=51235 $Y=56885
X3595 258 263 366 387 26 33 77 33 FA_X1 $T=56670 59800 0 180 $X=53515 $Y=58285
X3596 120 285 289 329 26 33 121 33 FA_X1 $T=54010 62600 1 0 $X=53895 $Y=61085
X3597 387 262 331 405 26 33 404 33 FA_X1 $T=54390 54200 1 0 $X=54275 $Y=52685
X3598 366 388 330 367 26 33 182 33 FA_X1 $T=54390 57000 0 0 $X=54275 $Y=56885
X3599 263 156 214 290 26 33 185 33 FA_X1 $T=56290 59800 0 0 $X=56175 $Y=59685
X3600 98 404 287 389 26 33 186 33 FA_X1 $T=56670 57000 1 0 $X=56555 $Y=55485
X3601 389 340 369 208 26 33 88 33 FA_X1 $T=58760 54200 1 0 $X=58645 $Y=52685
X3602 145 29 122 144 26 33 334 33 FA_X1 $T=58950 51400 0 0 $X=58835 $Y=51285
X3603 201 264 291 390 26 33 80 33 FA_X1 $T=61990 59800 0 180 $X=58835 $Y=58285
X3604 291 368 292 333 26 33 84 33 FA_X1 $T=59140 57000 0 0 $X=59025 $Y=56885
X3605 82 332 157 158 26 33 219 33 FA_X1 $T=59330 62600 1 0 $X=59215 $Y=61085
X3606 369 335 370 338 26 33 270 33 FA_X1 $T=61800 54200 1 0 $X=61685 $Y=52685
X3607 390 265 294 339 26 33 293 33 FA_X1 $T=62370 57000 1 0 $X=62255 $Y=55485
X3608 264 266 337 336 26 33 147 33 FA_X1 $T=62370 59800 0 0 $X=62255 $Y=59685
X3609 123 267 148 81 26 33 413 33 FA_X1 $T=62940 62600 1 0 $X=62825 $Y=61085
X3610 125 293 26 343 26 33 89 33 FA_X1 $T=64270 57000 0 0 $X=64155 $Y=56885
X3611 194 159 160 210 26 33 295 33 FA_X1 $T=65220 51400 0 0 $X=65105 $Y=51285
X3612 202 268 371 391 26 33 342 33 FA_X1 $T=65410 59800 0 0 $X=65295 $Y=59685
X3613 340 341 407 296 26 33 392 33 FA_X1 $T=66550 54200 0 0 $X=66435 $Y=54085
X3614 406 269 411 419 26 33 274 33 FA_X1 $T=68260 57000 1 0 $X=68145 $Y=55485
X3615 188 161 342 392 26 33 347 33 FA_X1 $T=71490 59800 1 180 $X=68335 $Y=59685
X3616 343 406 393 300 26 33 372 33 FA_X1 $T=69210 59800 1 0 $X=69095 $Y=58285
X3617 187 270 91 297 26 33 275 33 FA_X1 $T=69590 54200 0 0 $X=69475 $Y=54085
X3618 393 271 298 408 26 33 374 33 FA_X1 $T=71110 57000 0 0 $X=70995 $Y=56885
X3619 127 372 92 413 26 33 273 33 FA_X1 $T=71490 59800 0 0 $X=71375 $Y=59685
X3620 272 216 334 295 26 33 344 33 FA_X1 $T=72250 51400 0 0 $X=72135 $Y=51285
X3621 203 272 149 394 26 33 299 33 FA_X1 $T=72250 59800 1 0 $X=72135 $Y=58285
X3622 128 273 299 97 26 33 189 33 FA_X1 $T=74720 62600 1 0 $X=74605 $Y=61085
X3623 297 31 163 162 26 33 373 33 FA_X1 $T=75290 51400 0 0 $X=75175 $Y=51285
X3624 394 274 374 345 26 33 377 33 FA_X1 $T=75860 57000 1 0 $X=75745 $Y=55485
X3625 300 412 376 375 26 33 345 33 FA_X1 $T=81750 54200 0 180 $X=78595 $Y=52685
X3626 418 32 373 164 26 33 94 33 FA_X1 $T=78900 51400 0 0 $X=78785 $Y=51285
X3627 204 377 344 211 26 33 346 33 FA_X1 $T=78900 57000 1 0 $X=78785 $Y=55485
X3628 205 395 165 212 26 33 190 33 FA_X1 $T=78900 57000 0 0 $X=78785 $Y=56885
X3629 129 33 346 166 26 33 395 33 FA_X1 $T=84410 54200 1 180 $X=81255 $Y=54085
X3630 150 275 347 418 26 33 151 33 FA_X1 $T=81370 59800 0 0 $X=81255 $Y=59685
X3632 415 33 28 142 26 180 NAND3_X1 $T=42610 59800 0 0 $X=42495 $Y=59685
X3677 318 352 176 177 33 26 415 AND4_X1 $T=40900 54200 0 0 $X=40785 $Y=54085
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210
** N=440 EP=210 IP=5774 FDC=3090
M0 65 293 31 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=54195 $Y=50895 $D=1
M1 31 292 65 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54385 $Y=50895 $D=1
M2 31 290 291 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=54535 $Y=48690 $D=1
M3 65 246 31 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54575 $Y=50895 $D=1
M4 291 64 31 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54725 $Y=48690 $D=1
M5 31 246 65 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54765 $Y=50895 $D=1
M6 294 25 291 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54915 $Y=48690 $D=1
M7 65 292 31 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54955 $Y=50895 $D=1
M8 292 248 294 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=55105 $Y=48690 $D=1
M9 31 293 65 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=55145 $Y=50895 $D=1
M10 294 236 292 31 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=55295 $Y=48690 $D=1
M11 435 293 29 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=54195 $Y=50090 $D=0
M12 436 292 435 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54385 $Y=50090 $D=0
M13 437 290 29 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=54535 $Y=49280 $D=0
M14 65 246 436 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54575 $Y=50090 $D=0
M15 292 64 437 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54725 $Y=49280 $D=0
M16 438 246 65 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54765 $Y=50090 $D=0
M17 29 25 292 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54915 $Y=49280 $D=0
M18 439 292 438 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54955 $Y=50090 $D=0
M19 440 248 29 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=55105 $Y=49280 $D=0
M20 29 293 439 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=55145 $Y=50090 $D=0
M21 292 236 440 29 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=55295 $Y=49280 $D=0
X2686 366 224 31 29 282 OR2_X1 $T=35580 45800 0 0 $X=35465 $Y=45685
X2687 282 236 31 29 235 OR2_X1 $T=42990 48600 0 180 $X=42115 $Y=47085
X2688 64 242 31 29 236 OR2_X1 $T=52680 48600 1 180 $X=51805 $Y=48485
X2689 420 244 31 29 242 OR2_X1 $T=53250 45800 0 0 $X=53135 $Y=45685
X2741 403 10 31 29 20 DFF_X1 $T=1760 40200 0 0 $X=1645 $Y=40085
X2742 404 10 31 29 359 DFF_X1 $T=2330 43000 0 0 $X=2215 $Y=42885
X2743 407 11 31 29 86 DFF_X1 $T=2330 45800 1 0 $X=2215 $Y=44285
X2744 170 10 31 29 33 DFF_X1 $T=2520 51400 1 0 $X=2405 $Y=49885
X2745 218 11 31 29 113 DFF_X1 $T=3090 48600 0 0 $X=2975 $Y=48485
X2746 304 11 31 29 175 DFF_X1 $T=4610 48600 1 0 $X=4495 $Y=47085
X2747 405 10 31 29 305 DFF_X1 $T=5560 45800 1 0 $X=5445 $Y=44285
X2748 426 11 31 29 176 DFF_X1 $T=6320 48600 0 0 $X=6205 $Y=48485
X2749 171 10 31 29 221 DFF_X1 $T=6890 43000 1 0 $X=6775 $Y=41485
X2750 410 10 31 29 306 DFF_X1 $T=7840 43000 0 0 $X=7725 $Y=42885
X2751 358 10 31 29 301 DFF_X1 $T=7840 48600 1 0 $X=7725 $Y=47085
X2752 408 10 31 29 316 DFF_X1 $T=8790 45800 0 0 $X=8675 $Y=45685
X2753 172 10 31 29 114 DFF_X1 $T=14680 51400 1 0 $X=14565 $Y=49885
X2754 409 10 31 29 54 DFF_X1 $T=14870 45800 1 0 $X=14755 $Y=44285
X2755 406 10 31 29 219 DFF_X1 $T=15630 48600 0 0 $X=15515 $Y=48485
X2756 411 10 31 29 227 DFF_X1 $T=24940 48600 1 0 $X=24825 $Y=47085
X2757 220 11 31 29 93 DFF_X1 $T=25320 45800 0 0 $X=25205 $Y=45685
X2758 173 10 31 29 55 DFF_X1 $T=28550 51400 1 0 $X=28435 $Y=49885
X2788 34 1 31 29 403 31 AND2_X1 $T=1000 40200 0 0 $X=885 $Y=40085
X2789 32 4 31 29 426 31 AND2_X1 $T=1760 51400 0 180 $X=885 $Y=49885
X2790 34 2 31 29 404 31 AND2_X1 $T=1190 43000 1 0 $X=1075 $Y=41485
X2791 34 3 31 29 405 31 AND2_X1 $T=1190 45800 1 0 $X=1075 $Y=44285
X2792 32 5 31 29 407 31 AND2_X1 $T=1760 45800 0 0 $X=1645 $Y=45685
X2793 34 6 31 29 406 31 AND2_X1 $T=2520 51400 0 180 $X=1645 $Y=49885
X2794 34 9 31 29 408 31 AND2_X1 $T=3090 48600 0 180 $X=2215 $Y=47085
X2795 32 7 31 29 218 31 AND2_X1 $T=2330 48600 0 0 $X=2215 $Y=48485
X2796 32 8 31 29 304 31 AND2_X1 $T=2520 45800 0 0 $X=2405 $Y=45685
X2797 34 12 31 29 358 31 AND2_X1 $T=3850 48600 1 0 $X=3735 $Y=47085
X2798 34 13 31 29 409 31 AND2_X1 $T=4990 45800 0 0 $X=4875 $Y=45685
X2799 34 85 31 29 410 31 AND2_X1 $T=7080 43000 0 0 $X=6965 $Y=42885
X2800 32 14 31 29 220 31 AND2_X1 $T=8030 45800 0 0 $X=7915 $Y=45685
X2801 34 15 31 29 411 31 AND2_X1 $T=11830 48600 0 0 $X=11715 $Y=48485
X2802 372 226 31 29 228 31 AND2_X1 $T=36910 45800 0 180 $X=36035 $Y=44285
X2803 337 255 31 29 251 31 AND2_X1 $T=57810 45800 0 0 $X=57695 $Y=45685
X3141 318 21 367 222 31 29 OAI21_X1 $T=30260 43000 0 0 $X=30145 $Y=42885
X3142 121 22 368 56 31 29 OAI21_X1 $T=33680 45800 1 0 $X=33565 $Y=44285
X3143 414 223 370 369 31 29 OAI21_X1 $T=35010 48600 0 180 $X=34135 $Y=47085
X3144 325 228 232 327 31 29 OAI21_X1 $T=39000 48600 0 180 $X=38125 $Y=47085
X3145 281 282 234 248 31 29 OAI21_X1 $T=41090 48600 1 0 $X=40975 $Y=47085
X3146 287 241 416 243 31 29 OAI21_X1 $T=50400 48600 1 0 $X=50285 $Y=47085
X3147 288 242 123 290 31 29 OAI21_X1 $T=53630 48600 0 0 $X=53515 $Y=48485
X3148 338 253 341 340 31 29 OAI21_X1 $T=55530 48600 0 0 $X=55415 $Y=48485
X3149 66 251 256 342 31 29 OAI21_X1 $T=58950 48600 1 180 $X=58075 $Y=48485
X3252 322 31 29 223 31 INV_X1 $T=33870 45800 1 180 $X=33375 $Y=45685
X3253 321 31 29 369 31 INV_X1 $T=33870 48600 1 0 $X=33755 $Y=47085
X3254 368 31 29 281 31 INV_X1 $T=34820 45800 0 180 $X=34325 $Y=44285
X3255 370 31 29 325 31 INV_X1 $T=35010 48600 1 0 $X=34895 $Y=47085
X3256 278 31 29 327 31 INV_X1 $T=37100 48600 0 180 $X=36605 $Y=47085
X3257 415 31 29 328 31 INV_X1 $T=39570 45800 1 180 $X=39075 $Y=45685
X3258 234 31 29 288 31 INV_X1 $T=48690 48600 1 0 $X=48575 $Y=47085
X3259 289 31 29 253 31 INV_X1 $T=54580 45800 0 0 $X=54465 $Y=45685
X3260 252 31 29 340 31 INV_X1 $T=56100 45800 0 0 $X=55985 $Y=45685
X3261 341 31 29 66 31 INV_X1 $T=56290 48600 0 0 $X=56175 $Y=48485
X3262 343 31 29 342 31 INV_X1 $T=57810 48600 1 0 $X=57695 $Y=47085
X3263 344 31 29 380 31 INV_X1 $T=58570 45800 0 0 $X=58455 $Y=45685
X3472 318 202 203 31 29 277 31 HA_X1 $T=26080 43000 0 0 $X=25965 $Y=42885
X3473 323 324 190 31 29 372 31 HA_X1 $T=33870 43000 1 0 $X=33755 $Y=41485
X3474 226 191 329 31 29 280 31 HA_X1 $T=37480 43000 0 0 $X=37365 $Y=42885
X3475 230 284 60 31 29 241 31 HA_X1 $T=44890 45800 0 0 $X=44775 $Y=45685
X3544 20 37 31 29 INV_X2 $T=11260 40200 0 0 $X=11145 $Y=40085
X3545 221 47 31 29 INV_X2 $T=11830 40200 0 0 $X=11715 $Y=40085
X3546 86 87 31 29 INV_X2 $T=12020 45800 0 0 $X=11905 $Y=45685
X3547 359 42 31 29 INV_X2 $T=12210 43000 1 0 $X=12095 $Y=41485
X3548 113 36 31 29 INV_X2 $T=14870 48600 1 0 $X=14755 $Y=47085
X3549 175 38 31 29 INV_X2 $T=15440 48600 1 0 $X=15325 $Y=47085
X3550 219 26 31 29 INV_X2 $T=24370 48600 1 0 $X=24255 $Y=47085
X3551 305 57 31 29 INV_X2 $T=27410 45800 1 0 $X=27295 $Y=44285
X3552 301 53 31 29 INV_X2 $T=27980 48600 1 180 $X=27295 $Y=48485
X3553 114 84 31 29 INV_X2 $T=27980 51400 1 0 $X=27865 $Y=49885
X3554 306 43 31 29 INV_X2 $T=28550 43000 0 0 $X=28435 $Y=42885
X3555 316 79 31 29 INV_X2 $T=30070 45800 0 0 $X=29955 $Y=45685
X3556 227 61 31 29 INV_X2 $T=30260 48600 1 0 $X=30145 $Y=47085
X3557 54 28 31 29 INV_X2 $T=30640 45800 0 0 $X=30525 $Y=45685
X3558 55 78 31 29 INV_X2 $T=30640 48600 0 0 $X=30525 $Y=48485
X3656 29 414 133 395 31 31 XOR2_X1 $T=32730 48600 0 180 $X=31475 $Y=47085
X3657 29 281 164 367 31 31 XOR2_X1 $T=33110 45800 0 180 $X=31855 $Y=44285
X3658 29 325 94 373 31 31 XOR2_X1 $T=39380 48600 1 180 $X=38125 $Y=48485
X3659 29 288 122 416 31 31 XOR2_X1 $T=51920 48600 1 180 $X=50665 $Y=48485
X3660 29 338 102 339 31 31 XOR2_X1 $T=55720 51400 1 0 $X=55605 $Y=49885
X3668 318 31 21 222 29 31 NAND2_X1 $T=31400 45800 0 180 $X=30715 $Y=44285
X3669 323 31 277 322 29 31 NAND2_X1 $T=33680 45800 0 180 $X=32995 $Y=44285
X3670 287 31 241 243 29 31 NAND2_X1 $T=51730 48600 0 180 $X=51045 $Y=47085
X3671 379 31 302 289 29 31 NAND2_X1 $T=54010 45800 0 0 $X=53895 $Y=45685
X3672 58 29 37 307 31 31 NOR2_X1 $T=14300 43000 0 0 $X=14185 $Y=42885
X3673 36 29 185 161 31 31 NOR2_X1 $T=14680 40200 0 0 $X=14565 $Y=40085
X3674 87 29 40 39 31 31 NOR2_X1 $T=15250 40200 0 0 $X=15135 $Y=40085
X3675 41 29 42 308 31 31 NOR2_X1 $T=16010 43000 0 0 $X=15895 $Y=42885
X3676 38 29 43 268 31 31 NOR2_X1 $T=16580 40200 0 0 $X=16465 $Y=40085
X3677 116 29 57 360 31 31 NOR2_X1 $T=18100 45800 1 0 $X=17985 $Y=44285
X3678 80 29 49 310 31 31 NOR2_X1 $T=20000 45800 1 180 $X=19315 $Y=45685
X3679 44 29 47 46 31 31 NOR2_X1 $T=19810 40200 0 0 $X=19695 $Y=40085
X3680 45 29 79 271 31 31 NOR2_X1 $T=19810 45800 1 0 $X=19695 $Y=44285
X3681 44 29 48 311 31 31 NOR2_X1 $T=20000 45800 0 0 $X=19885 $Y=45685
X3682 107 29 28 362 31 31 NOR2_X1 $T=21330 45800 1 0 $X=21215 $Y=44285
X3683 80 29 48 272 31 31 NOR2_X1 $T=22280 45800 0 0 $X=22165 $Y=45685
X3684 35 29 50 273 31 31 NOR2_X1 $T=22850 45800 1 0 $X=22735 $Y=44285
X3685 36 29 49 274 31 31 NOR2_X1 $T=24750 45800 1 180 $X=24065 $Y=45685
X3686 44 29 52 275 31 31 NOR2_X1 $T=24750 51400 0 180 $X=24065 $Y=49885
X3687 68 29 53 427 31 31 NOR2_X1 $T=25320 45800 1 180 $X=24635 $Y=45685
X3688 17 29 18 313 31 31 NOR2_X1 $T=24750 51400 1 0 $X=24635 $Y=49885
X3689 91 29 77 364 31 31 NOR2_X1 $T=26080 43000 1 180 $X=25395 $Y=42885
X3690 17 29 47 163 31 31 NOR2_X1 $T=29120 40200 1 180 $X=28435 $Y=40085
X3691 318 29 21 366 31 31 NOR2_X1 $T=30260 45800 1 0 $X=30145 $Y=44285
X3692 17 29 185 319 31 31 NOR2_X1 $T=31780 40200 1 180 $X=31095 $Y=40085
X3693 44 29 40 320 31 31 NOR2_X1 $T=32350 40200 1 180 $X=31665 $Y=40085
X3694 87 29 52 147 31 31 NOR2_X1 $T=32350 51400 0 180 $X=31665 $Y=49885
X3695 223 29 321 395 31 31 NOR2_X1 $T=33490 45800 1 180 $X=32805 $Y=45685
X3696 323 29 277 321 31 31 NOR2_X1 $T=33680 43000 1 180 $X=32995 $Y=42885
X3697 17 29 78 326 31 31 NOR2_X1 $T=35770 51400 1 0 $X=35655 $Y=49885
X3698 44 29 76 371 31 31 NOR2_X1 $T=36910 51400 0 180 $X=36225 $Y=49885
X3699 226 29 372 278 31 31 NOR2_X1 $T=37480 45800 0 180 $X=36795 $Y=44285
X3700 17 29 40 279 31 31 NOR2_X1 $T=37100 40200 0 0 $X=36985 $Y=40085
X3701 228 29 278 373 31 31 NOR2_X1 $T=38240 48600 0 180 $X=37555 $Y=47085
X3702 230 29 280 415 31 31 NOR2_X1 $T=38430 45800 1 0 $X=38315 $Y=44285
X3703 44 29 37 231 31 31 NOR2_X1 $T=39380 43000 0 0 $X=39265 $Y=42885
X3704 36 29 97 149 31 31 NOR2_X1 $T=40520 51400 0 180 $X=39835 $Y=49885
X3705 80 29 59 178 31 31 NOR2_X1 $T=40520 51400 1 0 $X=40405 $Y=49885
X3706 56 29 235 246 31 31 NOR2_X1 $T=41090 45800 0 0 $X=40975 $Y=45685
X3707 36 29 43 330 31 31 NOR2_X1 $T=41850 43000 1 180 $X=41165 $Y=42885
X3708 36 29 84 237 31 31 NOR2_X1 $T=41470 51400 1 0 $X=41355 $Y=49885
X3709 87 29 57 238 31 31 NOR2_X1 $T=41660 45800 0 0 $X=41545 $Y=45685
X3710 80 29 42 331 31 31 NOR2_X1 $T=42610 40200 1 180 $X=41925 $Y=40085
X3711 58 29 79 376 31 31 NOR2_X1 $T=43750 45800 0 0 $X=43635 $Y=45685
X3712 87 29 59 398 31 31 NOR2_X1 $T=43940 48600 1 0 $X=43825 $Y=47085
X3713 41 29 28 428 31 31 NOR2_X1 $T=44320 45800 0 0 $X=44205 $Y=45685
X3714 58 29 97 283 31 31 NOR2_X1 $T=44320 48600 0 0 $X=44205 $Y=48485
X3715 17 29 61 285 31 31 NOR2_X1 $T=46030 48600 1 0 $X=45915 $Y=47085
X3716 44 29 78 334 31 31 NOR2_X1 $T=48500 48600 1 180 $X=47815 $Y=48485
X3717 80 29 76 378 31 31 NOR2_X1 $T=49070 48600 1 180 $X=48385 $Y=48485
X3718 17 29 77 336 31 31 NOR2_X1 $T=50210 48600 0 0 $X=50095 $Y=48485
X3719 287 29 241 244 31 31 NOR2_X1 $T=50970 45800 0 0 $X=50855 $Y=45685
X3720 379 29 302 252 31 31 NOR2_X1 $T=54390 45800 1 0 $X=54275 $Y=44285
X3721 253 29 252 339 31 31 NOR2_X1 $T=55530 45800 0 0 $X=55415 $Y=45685
X3722 17 29 37 153 31 31 NOR2_X1 $T=56290 40200 0 0 $X=56175 $Y=40085
X3723 255 29 337 343 31 31 NOR2_X1 $T=57240 45800 0 0 $X=57125 $Y=45685
X3724 251 29 343 103 31 31 NOR2_X1 $T=58190 48600 1 180 $X=57505 $Y=48485
X3725 247 29 249 344 31 31 NOR2_X1 $T=58190 48600 1 0 $X=58075 $Y=47085
X3726 44 29 42 104 31 31 NOR2_X1 $T=58950 40200 1 180 $X=58265 $Y=40085
X3727 80 29 43 126 31 31 NOR2_X1 $T=59140 43000 1 0 $X=59025 $Y=41485
X3728 73 29 48 181 31 31 NOR2_X1 $T=59900 51400 1 0 $X=59785 $Y=49885
X3729 41 29 50 258 31 31 NOR2_X1 $T=61420 43000 1 0 $X=61305 $Y=41485
X3730 17 29 28 296 31 31 NOR2_X1 $T=62370 48600 0 180 $X=61685 $Y=47085
X3731 44 29 28 382 31 31 NOR2_X1 $T=62940 45800 0 180 $X=62255 $Y=44285
X3732 17 29 79 346 31 31 NOR2_X1 $T=62370 45800 0 0 $X=62255 $Y=45685
X3733 71 29 49 105 31 31 NOR2_X1 $T=62940 51400 0 180 $X=62255 $Y=49885
X3734 38 29 53 432 31 31 NOR2_X1 $T=64270 43000 1 180 $X=63585 $Y=42885
X3735 68 29 26 383 31 31 NOR2_X1 $T=63700 48600 0 0 $X=63585 $Y=48485
X3736 116 29 77 297 31 31 NOR2_X1 $T=64460 43000 0 180 $X=63775 $Y=41485
X3737 36 29 57 384 31 31 NOR2_X1 $T=65030 43000 0 180 $X=64345 $Y=41485
X3738 91 29 18 402 31 31 NOR2_X1 $T=65030 48600 1 0 $X=64915 $Y=47085
X3739 58 29 28 385 31 31 NOR2_X1 $T=66170 43000 0 180 $X=65485 $Y=41485
X3740 71 29 48 387 31 31 NOR2_X1 $T=66550 45800 0 180 $X=65865 $Y=44285
X3741 73 29 52 388 31 31 NOR2_X1 $T=67880 45800 1 180 $X=67195 $Y=45685
X3742 35 29 26 69 31 31 NOR2_X1 $T=68070 51400 0 180 $X=67385 $Y=49885
X3743 17 29 43 349 31 31 NOR2_X1 $T=68830 43000 1 180 $X=68145 $Y=42885
X3744 45 29 84 262 31 31 NOR2_X1 $T=69210 45800 1 180 $X=68525 $Y=45685
X3745 35 29 97 351 31 31 NOR2_X1 $T=70350 48600 1 180 $X=69665 $Y=48485
X3746 68 29 18 129 31 31 NOR2_X1 $T=70350 51400 0 180 $X=69665 $Y=49885
X3747 17 29 42 299 31 31 NOR2_X1 $T=70160 43000 1 0 $X=70045 $Y=41485
X3748 107 29 59 352 31 31 NOR2_X1 $T=70350 48600 0 0 $X=70235 $Y=48485
X3749 91 29 52 75 31 31 NOR2_X1 $T=70350 51400 1 0 $X=70235 $Y=49885
X3750 17 29 57 265 31 31 NOR2_X1 $T=70540 45800 0 0 $X=70425 $Y=45685
X3751 116 29 76 390 31 31 NOR2_X1 $T=72440 48600 0 0 $X=72325 $Y=48485
X3752 41 29 61 354 31 31 NOR2_X1 $T=72440 51400 1 0 $X=72325 $Y=49885
X3753 38 29 78 392 31 31 NOR2_X1 $T=74530 48600 0 0 $X=74415 $Y=48485
X3754 44 29 57 168 31 31 NOR2_X1 $T=75670 40200 1 180 $X=74985 $Y=40085
X3755 44 29 79 391 31 31 NOR2_X1 $T=75290 48600 1 0 $X=75175 $Y=47085
X3756 80 29 79 130 31 31 NOR2_X1 $T=76430 43000 1 0 $X=76315 $Y=41485
X3757 36 29 50 355 31 31 NOR2_X1 $T=76620 48600 0 0 $X=76505 $Y=48485
X3758 80 29 28 393 31 31 NOR2_X1 $T=77000 45800 0 0 $X=76885 $Y=45685
X3759 87 29 53 356 31 31 NOR2_X1 $T=78140 48600 0 0 $X=78025 $Y=48485
X3760 58 29 77 394 31 31 NOR2_X1 $T=78140 51400 1 0 $X=78025 $Y=49885
X3761 281 222 414 366 31 29 31 AOI21_X1 $T=32920 45800 1 180 $X=32045 $Y=45685
X3762 322 222 229 224 31 29 31 AOI21_X1 $T=34820 45800 0 0 $X=34705 $Y=45685
X3763 230 280 375 415 31 29 31 AOI21_X1 $T=38430 45800 0 0 $X=38315 $Y=45685
X3764 288 243 338 244 31 29 31 AOI21_X1 $T=52300 48600 1 0 $X=52185 $Y=47085
X3765 289 243 250 420 31 29 31 AOI21_X1 $T=54200 48600 1 0 $X=54085 $Y=47085
X3766 247 249 431 344 31 29 31 AOI21_X1 $T=59520 48600 0 180 $X=58645 $Y=47085
X3767 24 29 359 306 31 315 31 NOR3_X1 $T=26840 43000 1 0 $X=26725 $Y=41485
X3768 22 29 121 235 31 293 31 NOR3_X1 $T=39950 45800 1 0 $X=39835 $Y=44285
X3769 31 375 179 232 29 31 XNOR2_X1 $T=40710 48600 0 0 $X=40595 $Y=48485
X3770 31 431 67 256 29 31 XNOR2_X1 $T=59900 51400 0 180 $X=58645 $Y=49885
X3773 114 29 219 118 33 363 31 31 NOR4_X1 $T=21900 51400 0 180 $X=20835 $Y=49885
X3774 221 29 19 20 305 276 31 31 NOR4_X1 $T=26080 40200 0 0 $X=25965 $Y=40085
X3775 316 29 301 227 55 317 31 31 NOR4_X1 $T=28930 48600 0 0 $X=28815 $Y=48485
X3776 88 307 308 268 29 31 309 31 FA_X1 $T=15820 43000 1 0 $X=15705 $Y=41485
X3777 115 16 269 118 29 31 143 31 FA_X1 $T=17910 51400 1 0 $X=17795 $Y=49885
X3778 269 311 310 113 29 31 412 31 FA_X1 $T=18290 48600 1 0 $X=18175 $Y=47085
X3779 89 314 270 309 29 31 144 31 FA_X1 $T=18860 43000 1 0 $X=18745 $Y=41485
X3780 117 412 132 361 29 31 119 31 FA_X1 $T=18860 48600 0 0 $X=18745 $Y=48485
X3781 312 360 271 362 29 31 270 31 FA_X1 $T=22470 43000 1 180 $X=19315 $Y=42885
X3782 361 272 274 86 29 31 120 31 FA_X1 $T=21330 48600 1 0 $X=21215 $Y=47085
X3783 162 51 413 312 29 31 145 31 FA_X1 $T=25320 43000 0 180 $X=22165 $Y=41485
X3784 90 219 313 275 29 31 30 31 FA_X1 $T=22280 48600 0 0 $X=22165 $Y=48485
X3785 413 273 427 364 29 31 314 31 FA_X1 $T=22470 43000 0 0 $X=22355 $Y=42885
X3786 225 221 319 320 29 31 174 31 FA_X1 $T=27600 43000 1 0 $X=27485 $Y=41485
X3787 329 23 207 134 29 31 324 31 FA_X1 $T=37100 40200 1 180 $X=33945 $Y=40085
X3788 177 227 326 371 29 31 148 31 FA_X1 $T=38240 48600 1 180 $X=35085 $Y=48485
X3789 165 225 24 279 29 31 374 31 FA_X1 $T=35770 43000 1 0 $X=35655 $Y=41485
X3790 396 231 331 330 29 31 31 31 FA_X1 $T=38810 43000 1 0 $X=38695 $Y=41485
X3791 95 233 396 19 29 31 208 31 FA_X1 $T=42040 40200 1 180 $X=38885 $Y=40085
X3792 150 237 398 283 29 31 239 31 FA_X1 $T=42040 51400 1 0 $X=41925 $Y=49885
X3793 166 397 31 374 29 31 377 31 FA_X1 $T=42230 43000 1 0 $X=42115 $Y=41485
X3794 240 209 96 135 29 31 284 31 FA_X1 $T=42230 43000 0 0 $X=42115 $Y=42885
X3795 233 238 376 428 29 31 397 31 FA_X1 $T=42230 45800 1 0 $X=42115 $Y=44285
X3796 332 204 98 377 29 31 151 31 FA_X1 $T=42610 40200 0 0 $X=42495 $Y=40085
X3797 99 285 334 378 29 31 399 31 FA_X1 $T=44890 48600 0 0 $X=44775 $Y=48485
X3798 180 239 399 335 29 31 100 31 FA_X1 $T=45080 51400 1 0 $X=44965 $Y=49885
X3799 333 136 63 419 29 31 400 31 FA_X1 $T=45270 43000 0 0 $X=45155 $Y=42885
X3800 245 192 332 206 29 31 286 31 FA_X1 $T=45650 40200 0 0 $X=45535 $Y=40085
X3801 302 240 400 286 29 31 287 31 FA_X1 $T=46790 45800 0 0 $X=46675 $Y=45685
X3802 335 193 301 336 29 31 152 31 FA_X1 $T=48120 51400 1 0 $X=48005 $Y=49885
X3803 254 137 62 417 29 31 401 31 FA_X1 $T=50020 43000 1 0 $X=49905 $Y=41485
X3804 337 418 333 401 29 31 379 31 FA_X1 $T=51350 45800 1 0 $X=51235 $Y=44285
X3805 430 245 124 139 29 31 418 31 FA_X1 $T=53060 43000 1 0 $X=52945 $Y=41485
X3806 417 138 101 194 29 31 419 31 FA_X1 $T=53250 40200 0 0 $X=53135 $Y=40085
X3807 295 254 125 186 29 31 257 31 FA_X1 $T=56100 43000 1 0 $X=55985 $Y=41485
X3808 167 303 345 195 29 31 154 31 FA_X1 $T=58950 40200 0 0 $X=58835 $Y=40085
X3809 249 257 430 196 29 31 255 31 FA_X1 $T=58950 45800 1 0 $X=58835 $Y=44285
X3810 381 305 346 382 29 31 261 31 FA_X1 $T=58950 45800 0 0 $X=58835 $Y=45685
X3811 29 381 316 296 29 31 127 31 FA_X1 $T=58950 48600 0 0 $X=58835 $Y=48485
X3812 303 258 432 297 29 31 128 31 FA_X1 $T=60660 43000 0 0 $X=60545 $Y=42885
X3813 345 384 197 385 29 31 155 31 FA_X1 $T=62370 40200 0 0 $X=62255 $Y=40085
X3814 347 387 199 93 29 31 386 31 FA_X1 $T=62940 45800 1 0 $X=62825 $Y=44285
X3815 259 347 298 429 29 31 205 31 FA_X1 $T=62940 45800 0 0 $X=62825 $Y=45685
X3816 182 259 198 140 29 31 156 31 FA_X1 $T=62940 51400 1 0 $X=62825 $Y=49885
X3817 433 260 359 349 29 31 72 31 FA_X1 $T=64270 43000 0 0 $X=64155 $Y=42885
X3818 298 383 402 388 29 31 264 31 FA_X1 $T=64270 48600 0 0 $X=64155 $Y=48485
X3819 260 20 299 187 29 31 157 31 FA_X1 $T=65410 40200 0 0 $X=65295 $Y=40085
X3820 429 262 352 351 29 31 389 31 FA_X1 $T=65600 48600 1 0 $X=65485 $Y=47085
X3821 70 261 348 74 29 31 357 31 FA_X1 $T=66550 45800 1 0 $X=66435 $Y=44285
X3822 348 27 108 306 29 31 421 31 FA_X1 $T=68450 40200 0 0 $X=68335 $Y=40085
X3823 158 421 106 386 29 31 350 31 FA_X1 $T=71870 43000 1 180 $X=68715 $Y=42885
X3824 353 263 141 210 29 31 422 31 FA_X1 $T=70730 43000 1 0 $X=70615 $Y=41485
X3825 183 264 389 300 29 31 263 31 FA_X1 $T=72250 48600 1 0 $X=72135 $Y=47085
X3826 109 160 295 423 29 31 247 31 FA_X1 $T=73960 45800 0 0 $X=73845 $Y=45685
X3827 131 354 392 390 29 31 300 31 FA_X1 $T=78140 51400 0 180 $X=74985 $Y=49885
X3828 31 422 81 350 29 31 423 31 FA_X1 $T=75860 43000 0 0 $X=75745 $Y=42885
X3829 82 265 391 393 29 31 267 31 FA_X1 $T=78710 48600 1 0 $X=78595 $Y=47085
X3830 112 355 356 394 29 31 266 31 FA_X1 $T=81750 48600 1 180 $X=78595 $Y=48485
X3831 110 200 111 424 29 31 31 31 FA_X1 $T=78900 43000 0 0 $X=78785 $Y=42885
X3832 434 266 267 433 29 31 424 31 FA_X1 $T=78900 45800 1 0 $X=78785 $Y=44285
X3833 169 201 31 188 29 31 160 31 FA_X1 $T=81370 40200 0 0 $X=81255 $Y=40085
X3834 83 29 357 434 29 31 425 31 FA_X1 $T=81370 45800 0 0 $X=81255 $Y=45685
X3835 184 425 353 142 29 31 159 31 FA_X1 $T=84410 51400 0 180 $X=81255 $Y=49885
X3838 365 31 315 92 29 189 NAND3_X1 $T=27220 51400 1 0 $X=27105 $Y=49885
X3839 369 31 327 328 29 224 NAND3_X1 $T=35960 48600 1 0 $X=35845 $Y=47085
X3840 340 31 342 380 29 420 NAND3_X1 $T=56860 48600 0 180 $X=55985 $Y=47085
X3842 230 280 29 229 228 31 328 248 AOI221_X1 $T=38430 45800 1 180 $X=37175 $Y=45685
X3843 247 249 29 250 251 31 380 290 AOI221_X1 $T=54960 48600 1 0 $X=54845 $Y=47085
X3851 363 146 317 276 31 29 365 AND4_X1 $T=25320 51400 1 0 $X=25205 $Y=49885
.ENDS
***************************************
.SUBCKT ICV_18 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 20 21
+ 22 23 24 25 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182
+ 183 184 185 186 187 188 189 190 191 192
** N=389 EP=190 IP=4512 FDC=2766
X2211 264 3 20 21 104 DFF_X1 $T=4610 40200 1 0 $X=4495 $Y=38685
X2212 310 3 20 21 157 DFF_X1 $T=7840 40200 1 0 $X=7725 $Y=38685
X2213 248 7 20 21 290 DFF_X1 $T=37860 31800 0 0 $X=37745 $Y=31685
X2246 22 89 20 21 264 20 AND2_X1 $T=1950 37400 1 180 $X=1075 $Y=37285
X2247 22 1 20 21 310 20 AND2_X1 $T=3090 40200 0 180 $X=2215 $Y=38685
X2248 22 2 20 21 103 20 AND2_X1 $T=3850 40200 1 0 $X=3735 $Y=38685
X2249 90 4 20 21 248 20 AND2_X1 $T=8410 37400 0 0 $X=8295 $Y=37285
X2831 104 48 20 21 INV_X2 $T=11070 40200 1 0 $X=10955 $Y=38685
X2832 157 27 20 21 INV_X2 $T=11640 40200 1 0 $X=11525 $Y=38685
X2833 54 99 20 21 INV_X2 $T=36150 31800 1 0 $X=36035 $Y=30285
X2834 88 13 20 21 INV_X2 $T=58380 31800 1 0 $X=58265 $Y=30285
X2835 290 70 20 21 INV_X2 $T=58950 31800 1 0 $X=58835 $Y=30285
X2921 23 21 48 311 20 20 NOR2_X1 $T=2330 37400 1 0 $X=2215 $Y=35885
X2922 24 21 51 265 20 20 NOR2_X1 $T=5940 34600 1 180 $X=5255 $Y=34485
X2923 25 21 30 339 20 20 NOR2_X1 $T=5940 37400 1 180 $X=5255 $Y=37285
X2924 82 21 27 314 20 20 NOR2_X1 $T=7840 34600 0 0 $X=7725 $Y=34485
X2925 28 21 29 313 20 20 NOR2_X1 $T=9930 34600 1 0 $X=9815 $Y=33085
X2926 98 21 37 211 20 20 NOR2_X1 $T=11640 37400 0 0 $X=11525 $Y=37285
X2927 33 21 12 212 20 20 NOR2_X1 $T=14110 31800 1 180 $X=13425 $Y=31685
X2928 31 21 32 268 20 20 NOR2_X1 $T=13920 37400 1 0 $X=13805 $Y=35885
X2929 33 21 34 316 20 20 NOR2_X1 $T=15060 34600 1 0 $X=14945 $Y=33085
X2930 79 21 12 317 20 20 NOR2_X1 $T=15820 37400 1 180 $X=15135 $Y=37285
X2931 35 21 39 318 20 20 NOR2_X1 $T=16960 31800 0 180 $X=16275 $Y=30285
X2932 91 21 39 364 20 20 NOR2_X1 $T=16580 37400 0 0 $X=16465 $Y=37285
X2933 36 21 29 214 20 20 NOR2_X1 $T=17530 40200 0 180 $X=16845 $Y=38685
X2934 35 21 44 341 20 20 NOR2_X1 $T=18860 34600 1 180 $X=18175 $Y=34485
X2935 45 21 40 384 20 20 NOR2_X1 $T=21330 31800 0 0 $X=21215 $Y=31685
X2936 41 21 43 273 20 20 NOR2_X1 $T=23040 31800 0 0 $X=22925 $Y=31685
X2937 13 21 47 274 20 20 NOR2_X1 $T=24940 31800 1 180 $X=24255 $Y=31685
X2938 45 21 43 217 20 20 NOR2_X1 $T=25130 37400 0 180 $X=24445 $Y=35885
X2939 119 21 46 114 20 20 NOR2_X1 $T=25890 31800 0 180 $X=25205 $Y=30285
X2940 41 21 47 275 20 20 NOR2_X1 $T=26460 34600 1 180 $X=25775 $Y=34485
X2941 13 21 78 276 20 20 NOR2_X1 $T=27220 37400 1 0 $X=27105 $Y=35885
X2942 36 21 27 277 20 20 NOR2_X1 $T=29120 37400 0 180 $X=28435 $Y=35885
X2943 28 21 48 278 20 20 NOR2_X1 $T=29690 34600 0 180 $X=29005 $Y=33085
X2944 126 21 27 279 20 20 NOR2_X1 $T=29500 40200 1 0 $X=29385 $Y=38685
X2945 119 21 72 325 20 20 NOR2_X1 $T=31210 31800 0 180 $X=30525 $Y=30285
X2946 70 21 46 326 20 20 NOR2_X1 $T=31210 31800 1 0 $X=31095 $Y=30285
X2947 82 21 51 280 20 20 NOR2_X1 $T=31970 34600 1 180 $X=31285 $Y=34485
X2948 36 21 51 221 20 20 NOR2_X1 $T=35010 37400 0 0 $X=34895 $Y=37285
X2949 28 21 30 289 20 20 NOR2_X1 $T=36720 34600 0 0 $X=36605 $Y=34485
X2950 82 21 37 380 20 20 NOR2_X1 $T=36910 37400 0 0 $X=36795 $Y=37285
X2951 33 21 43 230 20 20 NOR2_X1 $T=50970 31800 1 0 $X=50855 $Y=30285
X2952 119 21 74 120 20 20 NOR2_X1 $T=52110 31800 1 0 $X=51995 $Y=30285
X2953 91 21 47 349 20 20 NOR2_X1 $T=52680 31800 1 0 $X=52565 $Y=30285
X2954 35 21 78 332 20 20 NOR2_X1 $T=52870 34600 1 0 $X=52755 $Y=33085
X2955 23 21 32 233 20 20 NOR2_X1 $T=54770 31800 0 0 $X=54655 $Y=31685
X2956 98 21 39 234 20 20 NOR2_X1 $T=55530 37400 0 0 $X=55415 $Y=37285
X2957 31 21 44 334 20 20 NOR2_X1 $T=57050 37400 0 0 $X=56935 $Y=37285
X2958 24 21 12 294 20 20 NOR2_X1 $T=57240 34600 1 0 $X=57125 $Y=33085
X2959 25 21 34 387 20 20 NOR2_X1 $T=58380 31800 0 180 $X=57695 $Y=30285
X2960 41 21 67 263 20 20 NOR2_X1 $T=58380 31800 0 0 $X=58265 $Y=31685
X2961 79 21 40 376 20 20 NOR2_X1 $T=58950 37400 0 180 $X=58265 $Y=35885
X2962 13 21 75 297 20 20 NOR2_X1 $T=62940 31800 0 180 $X=62255 $Y=30285
X2963 99 21 74 382 20 20 NOR2_X1 $T=63510 31800 1 180 $X=62825 $Y=31685
X2964 31 21 43 237 20 20 NOR2_X1 $T=64080 37400 1 0 $X=63965 $Y=35885
X2965 91 21 71 335 20 20 NOR2_X1 $T=64650 34600 1 0 $X=64535 $Y=33085
X2966 82 21 12 100 20 20 NOR2_X1 $T=65600 40200 0 180 $X=64915 $Y=38685
X2967 79 21 47 300 20 20 NOR2_X1 $T=66740 34600 1 180 $X=66055 $Y=34485
X2968 33 21 78 256 20 20 NOR2_X1 $T=66930 37400 0 180 $X=66245 $Y=35885
X2969 45 21 72 255 20 20 NOR2_X1 $T=67120 34600 0 180 $X=66435 $Y=33085
X2970 13 21 73 149 20 20 NOR2_X1 $T=66550 37400 0 0 $X=66435 $Y=37285
X2971 35 21 46 301 20 20 NOR2_X1 $T=67690 31800 1 180 $X=67005 $Y=31685
X2972 35 21 67 353 20 20 NOR2_X1 $T=67690 34600 1 0 $X=67575 $Y=33085
X2973 45 21 75 388 20 20 NOR2_X1 $T=68260 34600 1 0 $X=68145 $Y=33085
X2974 126 21 37 150 20 20 NOR2_X1 $T=70350 40200 0 180 $X=69665 $Y=38685
X2975 41 21 74 355 20 20 NOR2_X1 $T=70730 34600 0 180 $X=70045 $Y=33085
X2976 25 21 43 389 20 20 NOR2_X1 $T=72250 34600 0 0 $X=72135 $Y=34485
X2977 31 21 78 336 20 20 NOR2_X1 $T=72250 40200 1 0 $X=72135 $Y=38685
X2978 98 21 47 378 20 20 NOR2_X1 $T=72630 37400 1 0 $X=72515 $Y=35885
X2979 82 21 39 240 20 20 NOR2_X1 $T=74340 37400 0 0 $X=74225 $Y=37285
X2980 23 21 44 305 20 20 NOR2_X1 $T=75290 34600 0 0 $X=75175 $Y=34485
X2981 24 21 40 337 20 20 NOR2_X1 $T=75480 37400 0 0 $X=75365 $Y=37285
X2982 28 21 34 304 20 20 NOR2_X1 $T=76620 37400 1 180 $X=75935 $Y=37285
X2983 28 21 12 83 20 20 NOR2_X1 $T=77760 31800 0 0 $X=77645 $Y=31685
X2984 168 21 290 54 20 18 20 NOR3_X1 $T=42610 31800 1 180 $X=41735 $Y=31685
X2986 358 359 312 170 21 20 137 20 FA_X1 $T=2330 31800 1 0 $X=2215 $Y=30285
X2987 340 122 313 314 21 20 312 20 FA_X1 $T=2330 34600 1 0 $X=2215 $Y=33085
X2988 244 311 265 339 21 20 359 20 FA_X1 $T=2330 34600 0 0 $X=2215 $Y=34485
X2989 266 360 340 245 21 20 210 20 FA_X1 $T=7460 37400 1 0 $X=7345 $Y=35885
X2990 245 184 315 123 21 20 105 20 FA_X1 $T=10310 31800 1 0 $X=10195 $Y=30285
X2991 246 210 358 362 21 20 344 20 FA_X1 $T=10500 31800 0 0 $X=10385 $Y=31685
X2992 269 213 267 244 21 20 247 20 FA_X1 $T=15250 34600 1 180 $X=12095 $Y=34485
X2993 267 211 268 317 21 20 361 20 FA_X1 $T=12210 37400 0 0 $X=12095 $Y=37285
X2994 315 212 106 318 21 20 107 20 FA_X1 $T=13350 31800 1 0 $X=13235 $Y=30285
X2995 319 214 171 124 21 20 360 20 FA_X1 $T=16960 40200 0 180 $X=13805 $Y=38685
X2996 362 342 270 361 21 20 138 20 FA_X1 $T=15250 31800 0 0 $X=15135 $Y=31685
X2997 213 316 364 341 21 20 270 20 FA_X1 $T=15250 34600 0 0 $X=15135 $Y=34485
X2998 363 365 266 38 21 20 271 20 FA_X1 $T=15820 37400 1 0 $X=15705 $Y=35885
X2999 365 247 322 185 21 20 366 20 FA_X1 $T=18290 31800 0 0 $X=18175 $Y=31685
X3000 343 215 108 172 21 20 109 20 FA_X1 $T=18860 31800 1 0 $X=18745 $Y=30285
X3001 383 366 344 165 21 20 110 20 FA_X1 $T=18860 34600 0 0 $X=18745 $Y=34485
X3002 111 216 383 343 21 20 218 20 FA_X1 $T=21900 37400 0 180 $X=18745 $Y=35885
X3003 284 20 271 246 21 20 321 20 FA_X1 $T=18860 37400 0 0 $X=18745 $Y=37285
X3004 320 125 319 173 21 20 272 20 FA_X1 $T=19050 40200 1 0 $X=18935 $Y=38685
X3005 379 384 273 274 21 20 342 20 FA_X1 $T=21330 34600 1 0 $X=21215 $Y=33085
X3006 158 218 321 166 21 20 139 20 FA_X1 $T=25130 40200 0 180 $X=21975 $Y=38685
X3007 112 190 113 379 21 20 322 20 FA_X1 $T=22280 31800 1 0 $X=22165 $Y=30285
X3008 42 217 275 276 21 20 367 20 FA_X1 $T=22280 34600 0 0 $X=22165 $Y=34485
X3009 346 219 272 167 21 20 20 20 FA_X1 $T=25320 37400 1 180 $X=22165 $Y=37285
X3010 219 5 345 367 21 20 215 20 FA_X1 $T=27410 34600 0 180 $X=24255 $Y=33085
X3011 323 324 115 279 21 20 220 20 FA_X1 $T=25130 40200 1 0 $X=25015 $Y=38685
X3012 347 220 320 174 21 20 368 20 FA_X1 $T=25320 37400 0 0 $X=25205 $Y=37285
X3013 140 6 326 325 21 20 345 20 FA_X1 $T=28930 31800 0 180 $X=25775 $Y=30285
X3014 324 277 278 280 21 20 369 20 FA_X1 $T=26460 34600 0 0 $X=26345 $Y=34485
X3015 222 175 346 368 21 20 281 20 FA_X1 $T=29120 37400 1 0 $X=29005 $Y=35885
X3016 370 127 369 269 21 20 285 20 FA_X1 $T=31780 31800 0 0 $X=31665 $Y=31685
X3017 282 49 284 281 21 20 50 20 FA_X1 $T=31970 37400 0 0 $X=31855 $Y=37285
X3018 283 370 177 176 21 20 288 20 FA_X1 $T=33110 31800 1 0 $X=32995 $Y=30285
X3019 291 286 288 363 21 20 92 20 FA_X1 $T=33680 34600 0 0 $X=33565 $Y=34485
X3020 286 285 93 52 21 20 216 20 FA_X1 $T=34820 31800 0 0 $X=34705 $Y=31685
X3021 287 221 289 380 21 20 224 20 FA_X1 $T=35580 37400 1 0 $X=35465 $Y=35885
X3022 226 222 327 254 21 20 223 20 FA_X1 $T=38620 37400 1 0 $X=38505 $Y=35885
X3023 385 8 178 283 21 20 371 20 FA_X1 $T=41850 31800 0 180 $X=38695 $Y=30285
X3024 94 223 291 371 21 20 225 20 FA_X1 $T=38810 34600 0 0 $X=38695 $Y=34485
X3025 160 225 282 250 21 20 53 20 FA_X1 $T=41850 37400 1 180 $X=38695 $Y=37285
X3026 249 224 116 323 21 20 327 20 FA_X1 $T=38810 40200 1 0 $X=38695 $Y=38685
X3027 159 226 385 331 21 20 142 20 FA_X1 $T=41660 37400 1 0 $X=41545 $Y=35885
X3028 95 179 347 128 21 20 372 20 FA_X1 $T=42230 31800 1 0 $X=42115 $Y=30285
X3029 227 56 55 191 21 20 329 20 FA_X1 $T=42230 34600 0 0 $X=42115 $Y=34485
X3030 141 57 96 328 21 20 58 20 FA_X1 $T=42230 37400 0 0 $X=42115 $Y=37285
X3031 328 9 97 372 21 20 250 20 FA_X1 $T=43180 31800 0 0 $X=43065 $Y=31685
X3032 373 129 117 333 21 20 251 20 FA_X1 $T=45270 31800 1 0 $X=45155 $Y=30285
X3033 306 227 251 330 21 20 60 20 FA_X1 $T=45270 34600 0 0 $X=45155 $Y=34485
X3034 59 61 156 329 21 20 143 20 FA_X1 $T=46790 34600 1 0 $X=46675 $Y=33085
X3035 330 228 118 386 21 20 252 20 FA_X1 $T=47930 40200 1 0 $X=47815 $Y=38685
X3036 295 229 252 62 21 20 144 20 FA_X1 $T=49450 37400 0 0 $X=49335 $Y=37285
X3037 229 63 348 65 21 20 331 20 FA_X1 $T=49830 34600 1 0 $X=49715 $Y=33085
X3038 155 230 349 332 21 20 231 20 FA_X1 $T=51730 31800 0 0 $X=51615 $Y=31685
X3039 386 232 292 287 21 20 348 20 FA_X1 $T=55340 37400 0 180 $X=52185 $Y=35885
X3040 161 10 249 374 21 20 145 20 FA_X1 $T=52490 37400 0 0 $X=52375 $Y=37285
X3041 374 231 293 375 21 20 254 20 FA_X1 $T=54010 34600 0 0 $X=53895 $Y=34485
X3042 333 186 180 130 21 20 253 20 FA_X1 $T=57810 31800 0 180 $X=54655 $Y=30285
X3043 292 233 294 387 21 20 375 20 FA_X1 $T=55340 31800 0 0 $X=55225 $Y=31685
X3044 232 234 334 376 21 20 293 20 FA_X1 $T=55340 37400 1 0 $X=55225 $Y=35885
X3045 162 11 121 169 21 20 228 20 FA_X1 $T=55720 40200 1 0 $X=55605 $Y=38685
X3046 351 253 298 350 21 20 64 20 FA_X1 $T=57810 34600 1 0 $X=57695 $Y=33085
X3047 352 263 297 382 21 20 298 20 FA_X1 $T=58950 31800 0 0 $X=58835 $Y=31685
X3048 377 235 351 131 21 20 236 20 FA_X1 $T=58950 37400 1 0 $X=58835 $Y=35885
X3049 69 236 295 68 21 20 66 20 FA_X1 $T=61990 37400 1 180 $X=58835 $Y=37285
X3050 296 352 299 381 21 20 147 20 FA_X1 $T=60850 34600 1 0 $X=60735 $Y=33085
X3051 381 237 300 256 21 20 238 20 FA_X1 $T=62370 34600 0 0 $X=62255 $Y=34485
X3052 235 238 181 132 21 20 148 20 FA_X1 $T=62370 37400 0 0 $X=62255 $Y=37285
X3053 146 187 188 290 21 20 239 20 FA_X1 $T=62940 31800 1 0 $X=62825 $Y=30285
X3054 299 335 301 255 21 20 350 20 FA_X1 $T=63510 31800 0 0 $X=63395 $Y=31685
X3055 242 133 192 296 21 20 257 20 FA_X1 $T=65600 40200 1 0 $X=65485 $Y=38685
X3056 356 134 14 15 21 20 258 20 FA_X1 $T=65980 31800 1 0 $X=65865 $Y=30285
X3057 354 353 388 355 21 20 303 20 FA_X1 $T=66740 34600 0 0 $X=66625 $Y=34485
X3058 163 354 356 259 21 20 76 20 FA_X1 $T=66930 37400 1 0 $X=66815 $Y=35885
X3059 302 239 303 258 21 20 260 20 FA_X1 $T=67690 31800 0 0 $X=67575 $Y=31685
X3060 77 260 182 377 21 20 241 20 FA_X1 $T=70730 34600 1 0 $X=70615 $Y=33085
X3061 259 389 378 336 21 20 357 20 FA_X1 $T=71300 37400 0 0 $X=71185 $Y=37285
X3062 151 135 136 304 21 20 261 20 FA_X1 $T=72820 40200 1 0 $X=72705 $Y=38685
X3063 81 16 189 373 21 20 262 20 FA_X1 $T=73390 31800 1 0 $X=73275 $Y=30285
X3064 80 240 305 337 21 20 338 20 FA_X1 $T=78900 34600 1 180 $X=75745 $Y=34485
X3065 164 257 307 183 21 20 243 20 FA_X1 $T=78330 31800 0 0 $X=78215 $Y=31685
X3066 101 241 86 262 21 20 152 20 FA_X1 $T=78900 34600 1 0 $X=78785 $Y=33085
X3067 85 243 306 309 21 20 84 20 FA_X1 $T=81940 34600 1 180 $X=78785 $Y=34485
X3068 21 242 308 302 21 20 153 20 FA_X1 $T=78900 40200 1 0 $X=78785 $Y=38685
X3069 307 17 102 87 21 20 154 20 FA_X1 $T=81370 31800 0 0 $X=81255 $Y=31685
X3070 308 357 338 261 21 20 309 20 FA_X1 $T=81370 37400 1 0 $X=81255 $Y=35885
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 30 31 32 33 34 36 37 38 39 41 42 43
+ 44 45 46 47 48 49 50 51 52 54 55 56 57 58 59 60 61 62 63 64
+ 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83 84
+ 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103 104
+ 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123 124
+ 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143 144
+ 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
** N=268 EP=156 IP=2841 FDC=1448
M0 47 45 11 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=54155 $Y=29090 $D=1
M1 11 7 47 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54345 $Y=29090 $D=1
M2 47 48 11 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54535 $Y=29090 $D=1
M3 11 46 47 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54725 $Y=29090 $D=1
M4 47 46 11 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=54915 $Y=29090 $D=1
M5 11 48 47 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=55105 $Y=29090 $D=1
M6 47 7 11 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=55295 $Y=29090 $D=1
M7 11 45 47 11 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=55485 $Y=29090 $D=1
M8 263 45 12 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=54155 $Y=29680 $D=0
M9 264 7 263 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54345 $Y=29680 $D=0
M10 265 48 264 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54535 $Y=29680 $D=0
M11 47 46 265 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54725 $Y=29680 $D=0
M12 266 46 47 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=54915 $Y=29680 $D=0
M13 267 48 266 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=55105 $Y=29680 $D=0
M14 268 7 267 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=55295 $Y=29680 $D=0
M15 12 45 268 12 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=55485 $Y=29680 $D=0
X1828 13 12 100 200 11 11 NOR2_X1 $T=2330 29000 1 0 $X=2215 $Y=27485
X1829 15 12 74 224 11 11 NOR2_X1 $T=5940 29000 0 180 $X=5255 $Y=27485
X1830 17 12 85 84 11 11 NOR2_X1 $T=8220 29000 1 0 $X=8105 $Y=27485
X1831 62 12 18 205 11 11 NOR2_X1 $T=9930 29000 0 0 $X=9815 $Y=28885
X1832 19 12 16 207 11 11 NOR2_X1 $T=13730 29000 0 180 $X=13045 $Y=27485
X1833 55 12 31 249 11 11 NOR2_X1 $T=14300 29000 0 180 $X=13615 $Y=27485
X1834 64 12 65 128 11 11 NOR2_X1 $T=15250 29000 0 0 $X=15135 $Y=28885
X1835 87 12 88 260 11 11 NOR2_X1 $T=17530 26200 1 0 $X=17415 $Y=24685
X1836 23 12 60 208 11 11 NOR2_X1 $T=19430 26200 1 180 $X=18745 $Y=26085
X1837 24 12 50 227 11 11 NOR2_X1 $T=20950 26200 1 180 $X=20265 $Y=26085
X1838 42 12 66 243 11 11 NOR2_X1 $T=24560 29000 1 180 $X=23875 $Y=28885
X1839 26 12 79 201 11 11 NOR2_X1 $T=25130 26200 0 180 $X=24445 $Y=24685
X1840 27 12 67 211 11 11 NOR2_X1 $T=26080 29000 1 0 $X=25965 $Y=27485
X1841 90 12 57 242 11 11 NOR2_X1 $T=26270 26200 1 0 $X=26155 $Y=24685
X1842 28 12 54 210 11 11 NOR2_X1 $T=27410 26200 0 180 $X=26725 $Y=24685
X1843 42 12 67 130 11 11 NOR2_X1 $T=27030 29000 0 0 $X=26915 $Y=28885
X1844 26 12 54 213 11 11 NOR2_X1 $T=28930 26200 1 180 $X=28245 $Y=26085
X1845 28 12 57 228 11 11 NOR2_X1 $T=28740 26200 1 0 $X=28625 $Y=24685
X1846 13 12 18 115 11 11 NOR2_X1 $T=29880 26200 0 180 $X=29195 $Y=24685
X1847 90 12 33 250 11 11 NOR2_X1 $T=31020 29000 0 180 $X=30335 $Y=27485
X1848 15 12 16 91 11 11 NOR2_X1 $T=31400 26200 0 180 $X=30715 $Y=24685
X1849 59 12 31 92 11 11 NOR2_X1 $T=32160 26200 1 0 $X=32045 $Y=24685
X1850 26 12 57 251 11 11 NOR2_X1 $T=33300 26200 0 180 $X=32615 $Y=24685
X1851 28 12 33 229 11 11 NOR2_X1 $T=33870 26200 0 180 $X=33185 $Y=24685
X1852 90 12 34 230 11 11 NOR2_X1 $T=33870 26200 1 0 $X=33755 $Y=24685
X1853 42 12 37 186 11 11 NOR2_X1 $T=36340 29000 0 0 $X=36225 $Y=28885
X1854 38 12 54 231 11 11 NOR2_X1 $T=38240 29000 0 0 $X=38125 $Y=28885
X1855 27 12 79 215 11 11 NOR2_X1 $T=39950 29000 0 180 $X=39265 $Y=27485
X1856 26 12 33 93 11 11 NOR2_X1 $T=40330 26200 0 180 $X=39645 $Y=24685
X1857 90 12 4 94 11 11 NOR2_X1 $T=40900 26200 0 0 $X=40785 $Y=26085
X1858 28 12 34 69 11 11 NOR2_X1 $T=42230 26200 1 0 $X=42115 $Y=24685
X1859 26 12 4 261 11 11 NOR2_X1 $T=42800 26200 1 0 $X=42685 $Y=24685
X1860 38 12 34 187 11 11 NOR2_X1 $T=43370 29000 1 0 $X=43255 $Y=27485
X1861 27 12 33 123 11 11 NOR2_X1 $T=44510 26200 0 0 $X=44395 $Y=26085
X1862 42 12 54 191 11 11 NOR2_X1 $T=50780 26200 0 0 $X=50665 $Y=26085
X1863 27 12 57 234 11 11 NOR2_X1 $T=51730 26200 1 0 $X=51615 $Y=24685
X1864 27 12 34 71 11 11 NOR2_X1 $T=55720 29000 0 0 $X=55605 $Y=28885
X1865 38 12 4 72 11 11 NOR2_X1 $T=56290 29000 0 0 $X=56175 $Y=28885
X1866 28 12 4 236 11 11 NOR2_X1 $T=57050 26200 0 180 $X=56365 $Y=24685
X1867 73 12 74 247 11 11 NOR2_X1 $T=58760 29000 0 0 $X=58645 $Y=28885
X1868 75 12 49 237 11 11 NOR2_X1 $T=59330 29000 0 0 $X=59215 $Y=28885
X1869 17 12 18 256 11 11 NOR2_X1 $T=61040 29000 0 180 $X=60355 $Y=27485
X1870 13 12 16 95 11 11 NOR2_X1 $T=61610 26200 0 180 $X=60925 $Y=24685
X1871 15 12 31 96 11 11 NOR2_X1 $T=63700 26200 0 180 $X=63015 $Y=24685
X1872 42 12 34 192 11 11 NOR2_X1 $T=63130 29000 1 0 $X=63015 $Y=27485
X1873 27 12 4 238 11 11 NOR2_X1 $T=65030 29000 1 0 $X=64915 $Y=27485
X1874 24 12 34 98 11 11 NOR2_X1 $T=65600 29000 1 180 $X=64915 $Y=28885
X1875 42 12 4 52 11 11 NOR2_X1 $T=67120 29000 1 180 $X=66435 $Y=28885
X1876 27 12 54 239 11 11 NOR2_X1 $T=67310 26200 0 180 $X=66625 $Y=24685
X1877 87 12 54 194 11 11 NOR2_X1 $T=67500 29000 1 0 $X=67385 $Y=27485
X1878 55 12 67 77 11 11 NOR2_X1 $T=68640 29000 1 180 $X=67955 $Y=28885
X1879 64 12 37 56 11 11 NOR2_X1 $T=70350 26200 0 180 $X=69665 $Y=24685
X1880 144 12 37 78 11 11 NOR2_X1 $T=70350 29000 1 180 $X=69665 $Y=28885
X1881 23 12 57 220 11 11 NOR2_X1 $T=70350 26200 1 0 $X=70235 $Y=24685
X1882 64 12 79 80 11 11 NOR2_X1 $T=70920 29000 1 180 $X=70235 $Y=28885
X1883 24 12 33 195 11 11 NOR2_X1 $T=72060 26200 1 180 $X=71375 $Y=26085
X1884 55 12 66 258 11 11 NOR2_X1 $T=71870 26200 1 0 $X=71755 $Y=24685
X1885 59 12 60 221 11 11 NOR2_X1 $T=74340 26200 0 0 $X=74225 $Y=26085
X1886 26 12 100 81 11 11 NOR2_X1 $T=75480 26200 1 0 $X=75365 $Y=24685
X1887 73 12 31 199 11 11 NOR2_X1 $T=76240 29000 0 0 $X=76125 $Y=28885
X1888 13 12 145 198 11 11 NOR2_X1 $T=77190 26200 1 0 $X=77075 $Y=24685
X1889 15 12 88 240 11 11 NOR2_X1 $T=77760 26200 0 0 $X=77645 $Y=26085
X1890 17 12 65 241 11 11 NOR2_X1 $T=78330 29000 0 0 $X=78215 $Y=28885
X1891 90 12 49 101 11 11 NOR2_X1 $T=78900 26200 1 0 $X=78785 $Y=24685
X1892 14 200 224 135 12 11 109 11 FA_X1 $T=2330 26200 1 0 $X=2215 $Y=24685
X1893 226 146 147 136 12 11 110 11 FA_X1 $T=2330 29000 0 0 $X=2215 $Y=28885
X1894 21 1 225 103 12 11 86 11 FA_X1 $T=8790 26200 0 0 $X=8675 $Y=26085
X1895 63 205 207 249 12 11 206 11 FA_X1 $T=10120 29000 1 0 $X=10005 $Y=27485
X1896 225 182 104 206 12 11 111 11 FA_X1 $T=17530 26200 0 180 $X=14375 $Y=24685
X1897 112 260 208 227 12 11 182 11 FA_X1 $T=18860 26200 1 180 $X=15705 $Y=26085
X1898 20 148 226 149 12 11 183 11 FA_X1 $T=15820 29000 1 0 $X=15705 $Y=27485
X1899 113 183 158 150 12 11 114 11 FA_X1 $T=18860 29000 1 0 $X=18745 $Y=27485
X1900 22 155 184 209 12 11 89 11 FA_X1 $T=20000 26200 1 0 $X=19885 $Y=24685
X1901 129 201 210 242 12 11 184 11 FA_X1 $T=22280 26200 0 0 $X=22165 $Y=26085
X1902 25 243 211 151 12 11 209 11 FA_X1 $T=22280 29000 1 0 $X=22165 $Y=27485
X1903 212 213 228 250 12 11 116 11 FA_X1 $T=26650 29000 1 0 $X=26535 $Y=27485
X1904 30 2 212 137 12 11 185 11 FA_X1 $T=30640 29000 1 180 $X=27485 $Y=28885
X1905 214 251 229 230 12 11 244 11 FA_X1 $T=28930 26200 0 0 $X=28815 $Y=26085
X1906 32 185 244 252 12 11 117 11 FA_X1 $T=33300 29000 0 0 $X=33185 $Y=28885
X1907 216 186 215 231 12 11 252 11 FA_X1 $T=36340 29000 1 0 $X=36225 $Y=27485
X1908 189 156 202 105 12 11 36 11 FA_X1 $T=39760 26200 0 180 $X=36605 $Y=24685
X1909 202 214 216 3 12 11 253 11 FA_X1 $T=37860 26200 0 0 $X=37745 $Y=26085
X1910 68 253 30 11 12 11 188 11 FA_X1 $T=38810 29000 0 0 $X=38695 $Y=28885
X1911 233 187 261 138 12 11 217 11 FA_X1 $T=41470 26200 0 0 $X=41355 $Y=26085
X1912 5 188 245 139 12 11 39 11 FA_X1 $T=42230 29000 0 0 $X=42115 $Y=28885
X1913 41 189 217 106 12 11 70 11 FA_X1 $T=46410 26200 0 180 $X=43255 $Y=24685
X1914 232 203 233 131 12 11 254 11 FA_X1 $T=43940 29000 1 0 $X=43825 $Y=27485
X1915 218 6 254 140 12 11 43 11 FA_X1 $T=49450 26200 0 180 $X=46295 $Y=24685
X1916 203 190 126 141 12 11 118 11 FA_X1 $T=50970 29000 0 0 $X=50855 $Y=28885
X1917 190 191 234 107 12 11 235 11 FA_X1 $T=51350 29000 1 0 $X=51235 $Y=27485
X1918 44 152 236 45 12 11 246 11 FA_X1 $T=53440 26200 1 0 $X=53325 $Y=24685
X1919 132 246 235 142 12 11 119 11 FA_X1 $T=57430 29000 0 180 $X=54275 $Y=27485
X1920 124 247 237 256 12 11 255 11 FA_X1 $T=57430 29000 1 0 $X=57315 $Y=27485
X1921 133 8 76 255 12 11 245 11 FA_X1 $T=58950 26200 0 0 $X=58835 $Y=26085
X1922 51 108 232 257 12 11 97 11 FA_X1 $T=61230 29000 0 0 $X=61115 $Y=28885
X1923 193 192 238 48 12 11 257 11 FA_X1 $T=62370 26200 0 0 $X=62255 $Y=26085
X1924 125 9 239 153 12 11 120 11 FA_X1 $T=63700 26200 1 0 $X=63585 $Y=24685
X1925 262 193 219 143 12 11 121 11 FA_X1 $T=65410 26200 0 0 $X=65295 $Y=26085
X1926 219 194 220 195 12 11 197 11 FA_X1 $T=68450 26200 0 0 $X=68335 $Y=26085
X1927 99 204 262 159 12 11 58 11 FA_X1 $T=70920 29000 0 0 $X=70805 $Y=28885
X1928 196 157 154 258 12 11 248 11 FA_X1 $T=75480 26200 0 180 $X=72325 $Y=24685
X1929 204 196 259 222 12 11 82 11 FA_X1 $T=75670 29000 1 0 $X=75555 $Y=27485
X1930 134 197 160 248 12 11 223 11 FA_X1 $T=78330 26200 0 0 $X=78215 $Y=26085
X1931 259 198 240 221 12 11 127 11 FA_X1 $T=78710 29000 1 0 $X=78595 $Y=27485
X1932 222 199 83 241 12 11 122 11 FA_X1 $T=78900 29000 0 0 $X=78785 $Y=28885
X1933 61 10 223 218 12 11 102 11 FA_X1 $T=84410 26200 1 180 $X=81255 $Y=26085
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 45 46 47 48 50 51 52 53 54 55 56 57 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
** N=281 EP=158 IP=3040 FDC=1590
M0 30 29 12 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=28885 $Y=22895 $D=1
M1 278 3 30 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29075 $Y=22895 $D=1
M2 12 177 278 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29265 $Y=22895 $D=1
M3 279 177 12 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29455 $Y=22895 $D=1
M4 30 3 279 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=29645 $Y=22895 $D=1
M5 12 29 30 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=6.225e-14 AS=5.81e-14 PD=1.13e-06 PS=1.11e-06 $X=29835 $Y=22895 $D=1
M6 280 179 12 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=6.225e-14 PD=1.11e-06 PS=1.13e-06 $X=30035 $Y=22895 $D=1
M7 30 180 280 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=30225 $Y=22895 $D=1
M8 281 180 30 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=30415 $Y=22895 $D=1
M9 12 179 281 12 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=30605 $Y=22895 $D=1
M10 198 29 199 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=28885 $Y=22090 $D=0
M11 13 3 198 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29075 $Y=22090 $D=0
M12 198 177 13 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29265 $Y=22090 $D=0
M13 13 177 198 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29455 $Y=22090 $D=0
M14 198 3 13 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=29645 $Y=22090 $D=0
M15 199 29 198 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=9.45e-14 AS=8.82e-14 PD=1.56e-06 PS=1.54e-06 $X=29835 $Y=22090 $D=0
M16 30 179 199 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=9.45e-14 PD=1.54e-06 PS=1.56e-06 $X=30035 $Y=22090 $D=0
M17 199 180 30 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=30225 $Y=22090 $D=0
M18 30 180 199 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=30415 $Y=22090 $D=0
M19 199 179 30 13 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=30605 $Y=22090 $D=0
X1410 68 4 12 13 94 OR2_X1 $T=32540 20600 1 0 $X=32425 $Y=19085
X1432 133 6 12 13 35 DFF_X1 $T=38620 20600 1 0 $X=38505 $Y=19085
X1433 88 174 12 13 179 12 AND2_X1 $T=21140 20600 0 180 $X=20265 $Y=19085
X1632 89 179 182 197 12 13 OAI21_X1 $T=28930 20600 1 0 $X=28815 $Y=19085
X1633 237 190 272 238 12 13 OAI21_X1 $T=71110 20600 0 0 $X=70995 $Y=20485
X1634 277 194 241 256 12 13 OAI21_X1 $T=82510 23400 0 180 $X=81635 $Y=21885
X1635 277 194 195 243 12 13 OAI21_X1 $T=84410 23400 1 180 $X=83535 $Y=23285
X1695 178 12 13 197 12 INV_X1 $T=27600 20600 1 0 $X=27485 $Y=19085
X1696 218 12 13 180 12 INV_X1 $T=29120 20600 0 0 $X=29005 $Y=20485
X1820 174 171 208 12 13 209 12 HA_X1 $T=14300 20600 0 0 $X=14185 $Y=20485
X1821 177 209 173 12 13 134 12 HA_X1 $T=16770 20600 0 0 $X=16655 $Y=20485
X1822 190 203 191 12 13 202 12 HA_X1 $T=72250 23400 1 0 $X=72135 $Y=21885
X1823 277 202 192 12 13 193 12 HA_X1 $T=77950 23400 1 0 $X=77835 $Y=21885
X1824 115 255 262 12 13 103 12 HA_X1 $T=81750 23400 0 180 $X=79735 $Y=21885
X1865 35 55 12 13 INV_X2 $T=42040 23400 1 0 $X=41925 $Y=21885
X1927 13 89 219 265 12 12 XOR2_X1 $T=30450 20600 1 0 $X=30335 $Y=19085
X1928 13 9 151 272 12 12 XOR2_X1 $T=70920 20600 1 0 $X=70805 $Y=19085
X1929 13 129 242 115 12 12 XOR2_X1 $T=82320 20600 1 0 $X=82205 $Y=19085
X1930 13 128 132 242 12 12 XOR2_X1 $T=84790 20600 0 180 $X=83535 $Y=19085
X1933 221 12 222 31 13 12 NAND2_X1 $T=33110 20600 0 0 $X=32995 $Y=20485
X1934 237 12 190 238 13 12 NAND2_X1 $T=71110 23400 1 0 $X=70995 $Y=21885
X1935 203 12 100 9 13 12 NAND2_X1 $T=74530 20600 0 180 $X=73845 $Y=19085
X1936 241 12 243 128 13 12 NAND2_X1 $T=82510 23400 1 0 $X=82395 $Y=21885
X1937 277 12 194 243 13 12 NAND2_X1 $T=83080 23400 0 0 $X=82965 $Y=23285
X1938 15 13 54 204 12 12 NOR2_X1 $T=5940 20600 1 180 $X=5255 $Y=20485
X1939 14 13 17 257 12 12 NOR2_X1 $T=6510 23400 1 0 $X=6395 $Y=21885
X1940 16 13 57 244 12 12 NOR2_X1 $T=7270 20600 1 180 $X=6585 $Y=20485
X1941 16 13 59 58 12 12 NOR2_X1 $T=7080 23400 0 0 $X=6965 $Y=23285
X1942 32 13 22 172 12 12 NOR2_X1 $T=16200 20600 0 0 $X=16085 $Y=20485
X1943 62 13 33 210 12 12 NOR2_X1 $T=19240 20600 1 180 $X=18555 $Y=20485
X1944 23 13 43 211 12 12 NOR2_X1 $T=19620 20600 0 180 $X=18935 $Y=19085
X1945 174 13 88 178 12 12 NOR2_X1 $T=21140 20600 1 0 $X=21025 $Y=19085
X1946 41 13 83 213 12 12 NOR2_X1 $T=22660 20600 1 0 $X=22545 $Y=19085
X1947 25 13 24 176 12 12 NOR2_X1 $T=24940 23400 0 180 $X=24255 $Y=21885
X1948 27 13 26 214 12 12 NOR2_X1 $T=25890 20600 1 180 $X=25205 $Y=20485
X1949 28 13 48 130 12 12 NOR2_X1 $T=25890 20600 0 0 $X=25775 $Y=20485
X1950 55 13 48 196 12 12 NOR2_X1 $T=26840 23400 0 180 $X=26155 $Y=21885
X1951 2 13 37 248 12 12 NOR2_X1 $T=27030 20600 1 180 $X=26345 $Y=20485
X1952 28 13 39 215 12 12 NOR2_X1 $T=26460 23400 0 0 $X=26345 $Y=23285
X1953 177 13 3 218 12 12 NOR2_X1 $T=26840 23400 1 0 $X=26725 $Y=21885
X1954 179 13 178 265 12 12 NOR2_X1 $T=27030 20600 0 0 $X=26915 $Y=20485
X1955 51 13 33 223 12 12 NOR2_X1 $T=34440 20600 1 0 $X=34325 $Y=19085
X1956 69 13 43 225 12 12 NOR2_X1 $T=36150 20600 0 0 $X=36035 $Y=20485
X1957 38 13 81 224 12 12 NOR2_X1 $T=36910 20600 1 0 $X=36795 $Y=19085
X1958 32 13 83 226 12 12 NOR2_X1 $T=39760 20600 0 0 $X=39645 $Y=20485
X1959 62 13 26 227 12 12 NOR2_X1 $T=40330 20600 0 0 $X=40215 $Y=20485
X1960 23 13 37 228 12 12 NOR2_X1 $T=42040 23400 0 180 $X=41355 $Y=21885
X1961 38 13 37 183 12 12 NOR2_X1 $T=43370 20600 1 180 $X=42685 $Y=20485
X1962 23 13 39 184 12 12 NOR2_X1 $T=43370 23400 1 0 $X=43255 $Y=21885
X1963 62 13 48 229 12 12 NOR2_X1 $T=44510 20600 0 0 $X=44395 $Y=20485
X1964 32 13 24 267 12 12 NOR2_X1 $T=45650 20600 1 180 $X=44965 $Y=20485
X1965 41 13 40 249 12 12 NOR2_X1 $T=46410 23400 0 180 $X=45725 $Y=21885
X1966 42 13 43 230 12 12 NOR2_X1 $T=51730 20600 0 0 $X=51615 $Y=20485
X1967 25 13 75 46 12 12 NOR2_X1 $T=54010 23400 0 0 $X=53895 $Y=23285
X1968 32 13 37 232 12 12 NOR2_X1 $T=54580 20600 1 0 $X=54465 $Y=19085
X1969 62 13 24 201 12 12 NOR2_X1 $T=55150 20600 1 0 $X=55035 $Y=19085
X1970 23 13 48 250 12 12 NOR2_X1 $T=55340 20600 0 0 $X=55225 $Y=20485
X1971 20 13 33 269 12 12 NOR2_X1 $T=61420 20600 0 180 $X=60735 $Y=19085
X1972 16 13 47 275 12 12 NOR2_X1 $T=61990 23400 0 180 $X=61305 $Y=21885
X1973 41 13 48 79 12 12 NOR2_X1 $T=64460 23400 0 0 $X=64345 $Y=23285
X1974 23 13 24 253 12 12 NOR2_X1 $T=66170 20600 0 180 $X=65485 $Y=19085
X1975 2 13 40 80 12 12 NOR2_X1 $T=67310 23400 1 180 $X=66625 $Y=23285
X1976 69 13 81 254 12 12 NOR2_X1 $T=69020 20600 1 180 $X=68335 $Y=20485
X1977 51 13 37 276 12 12 NOR2_X1 $T=68450 23400 1 0 $X=68335 $Y=21885
X1978 38 13 48 260 12 12 NOR2_X1 $T=69020 23400 1 0 $X=68905 $Y=21885
X1979 25 13 17 237 12 12 NOR2_X1 $T=70540 23400 1 0 $X=70425 $Y=21885
X1980 237 13 190 273 12 12 NOR2_X1 $T=71680 23400 1 0 $X=71565 $Y=21885
X1981 42 13 83 82 12 12 NOR2_X1 $T=72250 23400 0 0 $X=72135 $Y=23285
X1982 84 13 81 85 12 12 NOR2_X1 $T=72820 23400 0 0 $X=72705 $Y=23285
X1983 28 13 17 100 12 12 NOR2_X1 $T=73390 20600 1 0 $X=73275 $Y=19085
X1984 55 13 54 203 12 12 NOR2_X1 $T=73960 20600 0 0 $X=73845 $Y=20485
X1985 28 13 57 191 12 12 NOR2_X1 $T=74720 23400 0 180 $X=74035 $Y=21885
X1986 27 13 17 261 12 12 NOR2_X1 $T=75480 20600 0 180 $X=74795 $Y=19085
X1987 2 13 54 239 12 12 NOR2_X1 $T=76050 20600 0 180 $X=75365 $Y=19085
X1988 2 13 17 192 12 12 NOR2_X1 $T=75480 23400 1 0 $X=75365 $Y=21885
X1989 28 13 102 101 12 12 NOR2_X1 $T=77000 20600 1 0 $X=76885 $Y=19085
X1990 55 13 57 240 12 12 NOR2_X1 $T=77190 23400 0 0 $X=77075 $Y=23285
X1991 177 3 217 218 12 13 12 AOI21_X1 $T=28170 23400 0 180 $X=27295 $Y=21885
X1992 238 9 256 273 12 13 12 AOI21_X1 $T=71870 20600 0 0 $X=71755 $Y=20485
X1993 12 217 220 182 13 12 XNOR2_X1 $T=30830 23400 1 0 $X=30715 $Y=21885
X1994 12 256 136 195 13 12 XNOR2_X1 $T=83270 20600 0 0 $X=83155 $Y=20485
X1995 91 13 92 219 93 221 12 12 NOR4_X1 $T=31590 20600 1 0 $X=31475 $Y=19085
X1996 142 13 66 220 67 222 12 12 NOR4_X1 $T=31590 20600 0 0 $X=31475 $Y=20485
X1997 86 104 158 137 13 12 117 12 FA_X1 $T=2330 20600 1 0 $X=2215 $Y=19085
X1998 205 257 204 244 13 12 56 12 FA_X1 $T=2330 20600 0 0 $X=2215 $Y=20485
X1999 116 11 205 138 13 12 263 12 FA_X1 $T=2330 23400 0 0 $X=2215 $Y=23285
X2000 206 105 263 139 13 12 118 12 FA_X1 $T=5370 20600 1 0 $X=5255 $Y=19085
X2001 19 169 207 140 13 12 170 12 FA_X1 $T=9170 23400 0 0 $X=9055 $Y=23285
X2002 173 170 145 106 13 12 171 12 FA_X1 $T=9360 23400 1 0 $X=9245 $Y=21885
X2003 207 159 247 141 13 12 245 12 FA_X1 $T=12400 23400 1 0 $X=12285 $Y=21885
X2004 208 108 245 107 13 12 87 12 FA_X1 $T=12970 20600 1 0 $X=12855 $Y=19085
X2005 21 1 206 246 13 12 169 12 FA_X1 $T=15820 23400 0 0 $X=15705 $Y=23285
X2006 119 172 210 211 13 12 60 12 FA_X1 $T=16010 20600 1 0 $X=15895 $Y=19085
X2007 246 152 258 264 13 12 247 12 FA_X1 $T=18860 23400 1 0 $X=18745 $Y=21885
X2008 61 109 212 175 13 12 63 12 FA_X1 $T=18860 23400 0 0 $X=18745 $Y=23285
X2009 175 213 214 248 13 12 264 12 FA_X1 $T=22280 20600 0 0 $X=22165 $Y=20485
X2010 212 176 196 215 13 12 258 12 FA_X1 $T=22280 23400 0 0 $X=22165 $Y=23285
X2011 216 154 64 153 13 12 65 12 FA_X1 $T=27030 23400 0 0 $X=26915 $Y=23285
X2012 120 181 110 216 13 12 121 12 FA_X1 $T=30070 23400 0 0 $X=29955 $Y=23285
X2013 95 259 266 111 13 12 34 12 FA_X1 $T=35390 23400 1 0 $X=35275 $Y=21885
X2014 181 223 225 224 13 12 266 12 FA_X1 $T=39760 20600 1 180 $X=36605 $Y=20485
X2015 122 226 227 228 13 12 259 12 FA_X1 $T=38430 23400 1 0 $X=38315 $Y=21885
X2016 123 5 70 143 13 12 12 12 FA_X1 $T=38810 23400 0 0 $X=38695 $Y=23285
X2017 185 183 267 229 13 12 186 12 FA_X1 $T=42230 20600 1 0 $X=42115 $Y=19085
X2018 36 184 249 146 13 12 71 12 FA_X1 $T=42230 23400 0 0 $X=42115 $Y=23285
X2019 96 185 112 231 13 12 125 12 FA_X1 $T=45270 20600 1 0 $X=45155 $Y=19085
X2020 124 186 160 268 13 12 187 12 FA_X1 $T=45650 20600 0 0 $X=45535 $Y=20485
X2021 135 187 72 270 13 12 126 12 FA_X1 $T=47930 23400 0 0 $X=47815 $Y=23285
X2022 73 188 200 148 13 12 74 12 FA_X1 $T=50970 23400 0 0 $X=50855 $Y=23285
X2023 231 147 97 230 13 12 268 12 FA_X1 $T=54580 20600 0 180 $X=51425 $Y=19085
X2024 45 232 201 250 13 12 76 12 FA_X1 $T=58950 20600 1 180 $X=55795 $Y=20485
X2025 188 189 251 149 13 12 233 12 FA_X1 $T=55910 23400 0 0 $X=55795 $Y=23285
X2026 189 113 155 269 13 12 78 12 FA_X1 $T=57810 20600 1 0 $X=57695 $Y=19085
X2027 270 274 233 252 13 12 77 12 FA_X1 $T=61990 20600 1 180 $X=58835 $Y=20485
X2028 251 156 157 275 13 12 98 12 FA_X1 $T=58950 23400 0 0 $X=58835 $Y=23285
X2029 200 7 234 236 13 12 252 12 FA_X1 $T=65410 20600 1 180 $X=62255 $Y=20485
X2030 274 114 235 271 13 12 127 12 FA_X1 $T=62370 23400 1 0 $X=62255 $Y=21885
X2031 234 150 99 253 13 12 235 12 FA_X1 $T=62560 20600 1 0 $X=62445 $Y=19085
X2032 236 50 254 144 13 12 271 12 FA_X1 $T=65410 20600 0 0 $X=65295 $Y=20485
X2033 52 276 8 260 13 12 53 12 FA_X1 $T=67310 23400 0 0 $X=67195 $Y=23285
X2034 131 193 261 239 13 12 255 12 FA_X1 $T=78900 20600 0 0 $X=78785 $Y=20485
X2035 262 10 240 161 13 12 194 12 FA_X1 $T=78900 23400 0 0 $X=78785 $Y=23285
X2036 90 12 197 180 13 68 NAND3_X1 $T=29690 20600 1 0 $X=29575 $Y=19085
.ENDS
***************************************
.SUBCKT ICV_21
** N=2 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT ICV_22 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151
** N=257 EP=150 IP=3316 FDC=1490
X1551 182 7 16 17 47 DFF_X1 $T=38620 17800 1 0 $X=38505 $Y=16285
X1552 17 7 16 17 69 DFF_X1 $T=43180 17800 0 0 $X=43065 $Y=17685
X1553 226 7 16 17 50 DFF_X1 $T=52870 17800 1 0 $X=52755 $Y=16285
X1570 38 6 16 17 122 16 AND2_X1 $T=37860 17800 1 0 $X=37745 $Y=16285
X1571 38 60 16 17 182 16 AND2_X1 $T=40520 15000 1 180 $X=39645 $Y=14885
X1572 38 8 16 17 17 16 AND2_X1 $T=41090 15000 0 0 $X=40975 $Y=14885
X1573 38 9 16 17 226 16 AND2_X1 $T=44510 17800 1 0 $X=44395 $Y=16285
X1574 77 13 16 17 217 16 AND2_X1 $T=81560 17800 0 0 $X=81445 $Y=17685
X1763 188 162 200 64 16 17 OAI21_X1 $T=30070 17800 1 180 $X=29195 $Y=17685
X1764 65 163 240 161 16 17 OAI21_X1 $T=31400 15000 1 180 $X=30525 $Y=14885
X1765 211 173 212 56 16 17 OAI21_X1 $T=69590 17800 0 0 $X=69475 $Y=17685
X1766 105 14 249 103 16 17 OAI21_X1 $T=84410 15000 0 180 $X=83535 $Y=13485
X1824 221 16 17 162 16 INV_X1 $T=28740 17800 1 0 $X=28625 $Y=16285
X1825 200 16 17 139 16 INV_X1 $T=29310 17800 1 180 $X=28815 $Y=17685
X1826 222 16 17 64 16 INV_X1 $T=29690 17800 1 0 $X=29575 $Y=16285
X1827 47 16 17 4 16 INV_X1 $T=54200 17800 0 0 $X=54085 $Y=17685
X1828 50 16 17 48 16 INV_X1 $T=56100 17800 0 0 $X=55985 $Y=17685
X1829 212 16 17 215 16 INV_X1 $T=71300 17800 0 0 $X=71185 $Y=17685
X1922 181 149 256 16 17 24 16 HA_X1 $T=15630 17800 1 0 $X=15515 $Y=16285
X1923 105 112 176 16 17 101 16 HA_X1 $T=81940 15000 0 180 $X=79925 $Y=13485
X1960 69 28 16 17 INV_X2 $T=55530 17800 0 0 $X=55415 $Y=17685
X2019 17 188 33 247 16 16 XOR2_X1 $T=30070 17800 0 0 $X=29955 $Y=17685
X2020 17 5 84 240 16 16 XOR2_X1 $T=33490 17800 1 0 $X=33375 $Y=16285
X2021 17 78 218 249 16 16 XOR2_X1 $T=84790 15000 1 180 $X=83535 $Y=14885
X2023 181 16 31 221 17 16 NAND2_X1 $T=29310 15000 1 180 $X=28625 $Y=14885
X2024 65 16 163 161 17 16 NAND2_X1 $T=29310 15000 0 0 $X=29195 $Y=14885
X2025 68 17 52 235 16 16 NOR2_X1 $T=5940 15000 1 180 $X=5255 $Y=14885
X2026 39 17 18 189 16 16 NOR2_X1 $T=7270 15000 1 180 $X=6585 $Y=14885
X2027 19 17 49 190 16 16 NOR2_X1 $T=8600 15000 0 0 $X=8485 $Y=14885
X2028 45 17 20 191 16 16 NOR2_X1 $T=11830 17800 1 0 $X=11715 $Y=16285
X2029 21 17 41 178 16 16 NOR2_X1 $T=13920 17800 1 0 $X=13805 $Y=16285
X2030 23 17 36 245 16 16 NOR2_X1 $T=15630 15000 1 180 $X=14945 $Y=14885
X2031 40 17 62 192 16 16 NOR2_X1 $T=21710 15000 1 180 $X=21025 $Y=14885
X2032 40 17 42 239 16 16 NOR2_X1 $T=21330 17800 1 0 $X=21215 $Y=16285
X2033 55 17 3 194 16 16 NOR2_X1 $T=23420 17800 0 180 $X=22735 $Y=16285
X2034 55 17 42 220 16 16 NOR2_X1 $T=23040 15000 0 0 $X=22925 $Y=14885
X2035 48 17 27 238 16 16 NOR2_X1 $T=23420 17800 1 0 $X=23305 $Y=16285
X2036 48 17 3 246 16 16 NOR2_X1 $T=24180 15000 1 0 $X=24065 $Y=13485
X2037 28 17 3 151 16 16 NOR2_X1 $T=25320 15000 0 180 $X=24635 $Y=13485
X2038 30 17 27 128 16 16 NOR2_X1 $T=25320 15000 1 0 $X=25205 $Y=13485
X2039 28 17 27 160 16 16 NOR2_X1 $T=25890 17800 0 180 $X=25205 $Y=16285
X2040 4 17 29 81 16 16 NOR2_X1 $T=25890 15000 1 0 $X=25775 $Y=13485
X2041 28 17 29 198 16 16 NOR2_X1 $T=25890 17800 0 0 $X=25775 $Y=17685
X2042 30 17 29 199 16 16 NOR2_X1 $T=27030 17800 0 180 $X=26345 $Y=16285
X2043 30 17 63 196 16 16 NOR2_X1 $T=27030 17800 1 180 $X=26345 $Y=17685
X2044 4 17 63 180 16 16 NOR2_X1 $T=27600 17800 1 180 $X=26915 $Y=17685
X2045 28 17 42 82 16 16 NOR2_X1 $T=27790 15000 1 0 $X=27675 $Y=13485
X2046 181 17 31 222 16 16 NOR2_X1 $T=28170 15000 0 0 $X=28055 $Y=14885
X2047 162 17 222 247 16 16 NOR2_X1 $T=29120 17800 1 0 $X=29005 $Y=16285
X2048 30 17 3 32 16 16 NOR2_X1 $T=29310 15000 1 0 $X=29195 $Y=13485
X2049 4 17 27 83 16 16 NOR2_X1 $T=31020 15000 1 0 $X=30905 $Y=13485
X2050 65 17 163 34 16 16 NOR2_X1 $T=31400 15000 0 0 $X=31285 $Y=14885
X2051 40 17 36 164 16 16 NOR2_X1 $T=32730 15000 0 0 $X=32615 $Y=14885
X2052 55 17 10 201 16 16 NOR2_X1 $T=34630 15000 0 0 $X=34515 $Y=14885
X2053 68 17 41 223 16 16 NOR2_X1 $T=34630 17800 1 0 $X=34515 $Y=16285
X2054 48 17 37 202 16 16 NOR2_X1 $T=35200 15000 0 0 $X=35085 $Y=14885
X2055 19 17 10 257 16 16 NOR2_X1 $T=36910 17800 0 180 $X=36225 $Y=16285
X2056 28 17 62 165 16 16 NOR2_X1 $T=36910 15000 0 0 $X=36795 $Y=14885
X2057 39 17 36 203 16 16 NOR2_X1 $T=37860 17800 1 180 $X=37175 $Y=17685
X2058 30 17 42 224 16 16 NOR2_X1 $T=40520 15000 0 180 $X=39835 $Y=13485
X2059 4 17 3 225 16 16 NOR2_X1 $T=41090 15000 1 180 $X=40405 $Y=14885
X2060 40 17 41 166 16 16 NOR2_X1 $T=42800 15000 1 0 $X=42685 $Y=13485
X2061 55 17 36 183 16 16 NOR2_X1 $T=45080 15000 0 180 $X=44395 $Y=13485
X2062 48 17 10 204 16 16 NOR2_X1 $T=45840 15000 1 180 $X=45155 $Y=14885
X2063 28 17 37 167 16 16 NOR2_X1 $T=47170 15000 1 0 $X=47055 $Y=13485
X2064 19 17 42 205 16 16 NOR2_X1 $T=48120 17800 1 180 $X=47435 $Y=17685
X2065 4 17 42 184 16 16 NOR2_X1 $T=49830 15000 0 180 $X=49145 $Y=13485
X2066 45 17 3 227 16 16 NOR2_X1 $T=50020 17800 0 180 $X=49335 $Y=16285
X2067 21 17 27 241 16 16 NOR2_X1 $T=50210 17800 1 180 $X=49525 $Y=17685
X2068 28 17 10 168 16 16 NOR2_X1 $T=50970 15000 1 0 $X=50855 $Y=13485
X2069 46 17 10 67 16 16 NOR2_X1 $T=51730 17800 0 0 $X=51615 $Y=17685
X2070 68 17 37 88 16 16 NOR2_X1 $T=52300 17800 0 0 $X=52185 $Y=17685
X2071 30 17 37 242 16 16 NOR2_X1 $T=52680 15000 1 0 $X=52565 $Y=13485
X2072 4 17 62 206 16 16 NOR2_X1 $T=54580 15000 1 180 $X=53895 $Y=14885
X2073 48 17 36 89 16 16 NOR2_X1 $T=54580 15000 1 0 $X=54465 $Y=13485
X2074 40 17 49 90 16 16 NOR2_X1 $T=55150 15000 1 0 $X=55035 $Y=13485
X2075 28 17 36 207 16 16 NOR2_X1 $T=55720 15000 0 0 $X=55605 $Y=14885
X2076 30 17 10 208 16 16 NOR2_X1 $T=57620 15000 0 0 $X=57505 $Y=14885
X2077 68 17 36 71 16 16 NOR2_X1 $T=57810 17800 0 0 $X=57695 $Y=17685
X2078 4 17 37 209 16 16 NOR2_X1 $T=59710 17800 0 180 $X=59025 $Y=16285
X2079 39 17 10 92 16 16 NOR2_X1 $T=59330 17800 0 0 $X=59215 $Y=17685
X2080 51 17 52 228 16 16 NOR2_X1 $T=61420 17800 1 0 $X=61305 $Y=16285
X2081 35 17 11 185 16 16 NOR2_X1 $T=61990 17800 1 180 $X=61305 $Y=17685
X2082 44 17 12 229 16 16 NOR2_X1 $T=62940 15000 0 180 $X=62255 $Y=13485
X2083 35 17 27 93 16 16 NOR2_X1 $T=62370 17800 0 0 $X=62255 $Y=17685
X2084 40 17 18 248 16 16 NOR2_X1 $T=65980 17800 0 180 $X=65295 $Y=16285
X2085 44 17 29 95 16 16 NOR2_X1 $T=65980 17800 1 180 $X=65295 $Y=17685
X2086 55 17 49 186 16 16 NOR2_X1 $T=67120 15000 1 180 $X=66435 $Y=14885
X2087 48 17 20 250 16 16 NOR2_X1 $T=67310 17800 1 180 $X=66625 $Y=17685
X2088 45 17 62 96 16 16 NOR2_X1 $T=67310 17800 0 0 $X=67195 $Y=17685
X2089 23 17 3 97 16 16 NOR2_X1 $T=68450 17800 1 180 $X=67765 $Y=17685
X2090 35 17 72 98 16 16 NOR2_X1 $T=68070 15000 1 0 $X=67955 $Y=13485
X2091 28 17 20 210 16 16 NOR2_X1 $T=68830 15000 1 180 $X=68145 $Y=14885
X2092 30 17 72 211 16 16 NOR2_X1 $T=68450 17800 0 0 $X=68335 $Y=17685
X2093 4 17 11 173 16 16 NOR2_X1 $T=69020 17800 0 0 $X=68905 $Y=17685
X2094 44 17 11 127 16 16 NOR2_X1 $T=69970 15000 1 0 $X=69855 $Y=13485
X2095 30 17 41 213 16 16 NOR2_X1 $T=70540 15000 1 180 $X=69855 $Y=14885
X2096 51 17 12 73 16 16 NOR2_X1 $T=71110 15000 0 180 $X=70425 $Y=13485
X2097 4 17 36 172 16 16 NOR2_X1 $T=71110 15000 1 180 $X=70425 $Y=14885
X2098 40 17 72 231 16 16 NOR2_X1 $T=72820 17800 1 0 $X=72705 $Y=16285
X2099 51 17 72 232 16 16 NOR2_X1 $T=73010 15000 1 0 $X=72895 $Y=13485
X2100 55 17 11 233 16 16 NOR2_X1 $T=75100 17800 0 0 $X=74985 $Y=17685
X2101 48 17 12 252 16 16 NOR2_X1 $T=75670 17800 0 0 $X=75555 $Y=17685
X2102 28 17 52 253 16 16 NOR2_X1 $T=76240 15000 0 0 $X=76125 $Y=14885
X2103 28 17 12 175 16 16 NOR2_X1 $T=77570 17800 1 180 $X=76885 $Y=17685
X2104 30 17 18 234 16 16 NOR2_X1 $T=78330 17800 0 180 $X=77645 $Y=16285
X2105 30 17 52 216 16 16 NOR2_X1 $T=78330 17800 1 0 $X=78215 $Y=16285
X2106 4 17 49 255 16 16 NOR2_X1 $T=78710 15000 0 0 $X=78595 $Y=14885
X2107 221 161 129 138 16 17 16 AOI21_X1 $T=28170 17800 0 0 $X=28055 $Y=17685
X2108 161 5 188 34 16 17 16 AOI21_X1 $T=31780 17800 1 0 $X=31665 $Y=16285
X2109 58 17 215 74 16 214 16 NOR3_X1 $T=72440 17800 1 180 $X=71565 $Y=17685
X2110 79 217 16 78 77 13 17 OAI22_X1 $T=83270 17800 1 180 $X=82205 $Y=17685
X2111 143 17 104 218 102 187 16 16 NOR4_X1 $T=84410 17800 0 180 $X=83345 $Y=16285
X2112 15 235 189 190 17 16 113 16 FA_X1 $T=2330 15000 0 0 $X=2215 $Y=14885
X2113 134 106 107 141 17 16 157 16 FA_X1 $T=2330 17800 1 0 $X=2215 $Y=16285
X2114 135 157 236 144 17 16 114 16 FA_X1 $T=5750 17800 1 0 $X=5635 $Y=16285
X2115 115 193 80 244 17 16 243 16 FA_X1 $T=8790 17800 1 0 $X=8675 $Y=16285
X2116 236 1 243 108 17 16 219 16 FA_X1 $T=9740 15000 1 0 $X=9625 $Y=13485
X2117 136 158 61 237 17 16 116 16 FA_X1 $T=11640 17800 0 0 $X=11525 $Y=17685
X2118 237 191 178 245 17 16 244 16 FA_X1 $T=12020 15000 0 0 $X=11905 $Y=14885
X2119 256 2 219 145 17 16 163 16 FA_X1 $T=15820 15000 0 180 $X=12665 $Y=13485
X2120 25 159 146 197 17 16 117 16 FA_X1 $T=18860 15000 0 180 $X=15705 $Y=13485
X2121 26 147 195 179 17 16 159 16 FA_X1 $T=19620 15000 1 180 $X=16465 $Y=14885
X2122 179 192 220 246 17 16 118 16 FA_X1 $T=18860 15000 1 0 $X=18745 $Y=13485
X2123 158 239 194 238 17 16 193 16 FA_X1 $T=18860 17800 0 0 $X=18745 $Y=17685
X2124 137 198 196 150 17 16 197 16 FA_X1 $T=22280 17800 0 0 $X=22165 $Y=17685
X2125 195 160 199 180 17 16 119 16 FA_X1 $T=23610 15000 0 0 $X=23495 $Y=14885
X2126 120 164 201 202 17 16 121 16 FA_X1 $T=33870 15000 1 0 $X=33755 $Y=13485
X2127 140 223 203 257 17 16 85 16 FA_X1 $T=34250 17800 0 0 $X=34135 $Y=17685
X2128 130 165 224 225 17 16 123 16 FA_X1 $T=36910 15000 1 0 $X=36795 $Y=13485
X2129 131 166 183 204 17 16 86 16 FA_X1 $T=42230 15000 0 0 $X=42115 $Y=14885
X2130 87 205 227 241 17 16 124 16 FA_X1 $T=45270 17800 1 0 $X=45155 $Y=16285
X2131 66 167 148 184 17 16 133 16 FA_X1 $T=45840 15000 0 0 $X=45725 $Y=14885
X2132 43 168 242 206 17 16 125 16 FA_X1 $T=50970 15000 0 0 $X=50855 $Y=14885
X2133 70 207 208 209 17 16 126 16 FA_X1 $T=56100 17800 1 0 $X=55985 $Y=16285
X2134 91 169 110 109 17 16 17 16 FA_X1 $T=58950 15000 1 0 $X=58835 $Y=13485
X2135 169 185 229 228 17 16 171 16 FA_X1 $T=59710 15000 0 0 $X=59595 $Y=14885
X2136 53 248 186 250 17 16 170 16 FA_X1 $T=62370 17800 1 0 $X=62255 $Y=16285
X2137 94 170 171 230 17 16 54 16 FA_X1 $T=62940 15000 1 0 $X=62825 $Y=13485
X2138 230 210 213 172 17 16 57 16 FA_X1 $T=65980 17800 1 0 $X=65865 $Y=16285
X2139 76 174 251 232 17 16 59 16 FA_X1 $T=76240 15000 1 180 $X=73085 $Y=14885
X2140 251 231 233 252 17 16 177 16 FA_X1 $T=74720 17800 1 0 $X=74605 $Y=16285
X2141 174 253 234 255 17 16 176 16 FA_X1 $T=77000 15000 1 0 $X=76885 $Y=13485
X2142 254 175 216 142 17 16 77 16 FA_X1 $T=78520 17800 0 0 $X=78405 $Y=17685
X2143 132 177 111 254 17 16 14 16 FA_X1 $T=81940 17800 0 180 $X=78785 $Y=16285
X2145 187 16 214 99 100 75 17 NAND4_X1 $T=71870 17800 1 0 $X=71755 $Y=16285
.ENDS
***************************************
.SUBCKT ICV_23 1 2 3 4 5 6 7 8 9 10 11 12 13 15 16 17 18 19 20 21
+ 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145
** N=264 EP=144 IP=2924 FDC=1594
X1605 240 11 12 127 11 INV_X1 $T=83650 9400 0 180 $X=83155 $Y=7885
X1730 263 96 9 11 12 80 11 HA_X1 $T=81940 12200 0 180 $X=79925 $Y=10685
X1803 12 240 117 231 11 11 XOR2_X1 $T=84790 12200 0 180 $X=83535 $Y=10685
X1805 263 11 185 66 12 11 NAND2_X1 $T=80800 9400 1 0 $X=80685 $Y=7885
X1806 68 11 50 81 12 11 NAND2_X1 $T=82320 12200 0 0 $X=82205 $Y=12085
X1807 13 12 30 210 11 11 NOR2_X1 $T=5940 9400 0 180 $X=5255 $Y=7885
X1808 53 12 15 232 11 11 NOR2_X1 $T=6510 9400 0 0 $X=6395 $Y=9285
X1809 13 12 15 71 11 11 NOR2_X1 $T=8410 9400 1 0 $X=8295 $Y=7885
X1810 31 12 47 165 11 11 NOR2_X1 $T=10500 12200 1 0 $X=10385 $Y=10685
X1811 16 12 23 243 11 11 NOR2_X1 $T=12400 9400 0 0 $X=12285 $Y=9285
X1812 17 12 4 187 11 11 NOR2_X1 $T=13540 9400 1 180 $X=12855 $Y=9285
X1813 17 12 23 253 11 11 NOR2_X1 $T=13540 9400 0 0 $X=13425 $Y=9285
X1814 21 12 18 166 11 11 NOR2_X1 $T=15820 12200 0 0 $X=15705 $Y=12085
X1815 21 12 4 167 11 11 NOR2_X1 $T=17150 9400 0 0 $X=17035 $Y=9285
X1816 28 12 18 212 11 11 NOR2_X1 $T=18290 9400 1 180 $X=17605 $Y=9285
X1817 28 12 24 213 11 11 NOR2_X1 $T=18100 12200 1 0 $X=17985 $Y=10685
X1818 33 12 24 254 11 11 NOR2_X1 $T=18860 9400 1 180 $X=18175 $Y=9285
X1819 33 12 20 246 11 11 NOR2_X1 $T=18670 12200 1 0 $X=18555 $Y=10685
X1820 39 12 20 214 11 11 NOR2_X1 $T=21520 12200 0 180 $X=20835 $Y=10685
X1821 46 12 35 233 11 11 NOR2_X1 $T=22280 12200 0 0 $X=22165 $Y=12085
X1822 27 12 22 255 11 11 NOR2_X1 $T=24180 12200 1 180 $X=23495 $Y=12085
X1823 21 12 23 190 11 11 NOR2_X1 $T=24180 9400 1 0 $X=24065 $Y=7885
X1824 33 12 18 215 11 11 NOR2_X1 $T=26650 12200 0 180 $X=25965 $Y=10685
X1825 28 12 4 235 11 11 NOR2_X1 $T=26840 9400 0 180 $X=26155 $Y=7885
X1826 39 12 24 191 11 11 NOR2_X1 $T=28550 9400 0 0 $X=28435 $Y=9285
X1827 46 12 20 192 11 11 NOR2_X1 $T=31590 12200 0 180 $X=30905 $Y=10685
X1828 27 12 35 216 11 11 NOR2_X1 $T=32160 12200 0 180 $X=31475 $Y=10685
X1829 31 12 78 236 11 11 NOR2_X1 $T=32350 9400 0 0 $X=32235 $Y=9285
X1830 21 12 47 170 11 11 NOR2_X1 $T=33300 12200 0 0 $X=33185 $Y=12085
X1831 28 12 23 193 11 11 NOR2_X1 $T=34820 12200 1 0 $X=34705 $Y=10685
X1832 33 12 4 247 11 11 NOR2_X1 $T=37480 12200 1 180 $X=36795 $Y=12085
X1833 29 12 30 196 11 11 NOR2_X1 $T=37860 12200 1 0 $X=37745 $Y=10685
X1834 59 12 15 256 11 11 NOR2_X1 $T=38240 9400 0 0 $X=38125 $Y=9285
X1835 31 12 30 173 11 11 NOR2_X1 $T=40520 12200 0 180 $X=39835 $Y=10685
X1836 17 12 37 237 11 11 NOR2_X1 $T=41090 9400 1 0 $X=40975 $Y=7885
X1837 16 12 78 248 11 11 NOR2_X1 $T=42800 9400 1 180 $X=42115 $Y=9285
X1838 21 12 42 262 11 11 NOR2_X1 $T=44890 9400 0 180 $X=44205 $Y=7885
X1839 28 12 47 219 11 11 NOR2_X1 $T=46410 12200 1 180 $X=45725 $Y=12085
X1840 33 12 23 257 11 11 NOR2_X1 $T=46980 12200 1 180 $X=46295 $Y=12085
X1841 29 12 15 75 11 11 NOR2_X1 $T=48500 9400 0 180 $X=47815 $Y=7885
X1842 21 12 37 175 11 11 NOR2_X1 $T=48120 9400 0 0 $X=48005 $Y=9285
X1843 45 12 35 34 11 11 NOR2_X1 $T=49070 12200 1 180 $X=48385 $Y=12085
X1844 28 12 42 199 11 11 NOR2_X1 $T=49640 9400 0 0 $X=49525 $Y=9285
X1845 33 12 47 258 11 11 NOR2_X1 $T=51540 9400 1 180 $X=50855 $Y=9285
X1846 39 12 23 176 11 11 NOR2_X1 $T=51540 12200 1 0 $X=51425 $Y=10685
X1847 46 12 4 200 11 11 NOR2_X1 $T=52300 12200 0 0 $X=52185 $Y=12085
X1848 27 12 4 202 11 11 NOR2_X1 $T=56670 12200 0 0 $X=56555 $Y=12085
X1849 21 12 78 177 11 11 NOR2_X1 $T=57050 9400 0 0 $X=56935 $Y=9285
X1850 46 12 23 203 11 11 NOR2_X1 $T=57430 12200 1 0 $X=57315 $Y=10685
X1851 28 12 37 222 11 11 NOR2_X1 $T=58760 12200 1 0 $X=58645 $Y=10685
X1852 33 12 42 204 11 11 NOR2_X1 $T=59330 9400 1 0 $X=59215 $Y=7885
X1853 17 12 30 60 11 11 NOR2_X1 $T=60280 12200 0 0 $X=60165 $Y=12085
X1854 16 12 15 61 11 11 NOR2_X1 $T=60850 12200 0 0 $X=60735 $Y=12085
X1855 62 12 4 180 11 11 NOR2_X1 $T=63510 12200 0 0 $X=63395 $Y=12085
X1856 44 12 24 260 11 11 NOR2_X1 $T=66930 12200 1 180 $X=66245 $Y=12085
X1857 17 12 15 226 11 11 NOR2_X1 $T=67120 9400 0 180 $X=66435 $Y=7885
X1858 45 12 18 227 11 11 NOR2_X1 $T=67120 12200 0 180 $X=66435 $Y=10685
X1859 39 12 37 181 11 11 NOR2_X1 $T=68830 12200 1 0 $X=68715 $Y=10685
X1860 46 12 42 252 11 11 NOR2_X1 $T=70160 12200 1 0 $X=70045 $Y=10685
X1861 27 12 47 183 11 11 NOR2_X1 $T=71490 12200 1 0 $X=71375 $Y=10685
X1862 39 12 30 228 11 11 NOR2_X1 $T=72820 12200 1 180 $X=72135 $Y=12085
X1863 33 12 30 63 11 11 NOR2_X1 $T=72440 9400 1 0 $X=72325 $Y=7885
X1864 39 12 78 205 11 11 NOR2_X1 $T=72630 9400 0 0 $X=72515 $Y=9285
X1865 46 12 37 238 11 11 NOR2_X1 $T=74530 9400 0 0 $X=74415 $Y=9285
X1866 46 12 78 206 11 11 NOR2_X1 $T=74530 12200 1 0 $X=74415 $Y=10685
X1867 27 12 42 261 11 11 NOR2_X1 $T=75670 9400 1 180 $X=74985 $Y=9285
X1868 27 12 37 207 11 11 NOR2_X1 $T=75670 12200 0 180 $X=74985 $Y=10685
X1869 62 12 47 65 11 11 NOR2_X1 $T=76050 9400 1 0 $X=75935 $Y=7885
X1870 62 12 42 184 11 11 NOR2_X1 $T=77000 12200 0 0 $X=76885 $Y=12085
X1871 44 12 4 49 11 11 NOR2_X1 $T=77570 9400 1 0 $X=77455 $Y=7885
X1872 45 12 23 126 11 11 NOR2_X1 $T=77570 9400 0 0 $X=77455 $Y=9285
X1873 44 12 23 208 11 11 NOR2_X1 $T=77570 12200 0 0 $X=77455 $Y=12085
X1874 45 12 47 230 11 11 NOR2_X1 $T=79470 12200 1 180 $X=78785 $Y=12085
X1875 263 12 185 67 11 11 NOR2_X1 $T=81370 9400 1 0 $X=81255 $Y=7885
X1876 68 12 50 209 11 11 NOR2_X1 $T=83840 12200 0 0 $X=83725 $Y=12085
X1877 263 185 231 67 11 12 11 AOI21_X1 $T=81180 9400 0 0 $X=81065 $Y=9285
X1878 81 10 240 209 11 12 11 AOI21_X1 $T=83650 9400 0 0 $X=83535 $Y=9285
X1879 10 12 209 83 11 82 11 NOR3_X1 $T=84410 9400 0 180 $X=83535 $Y=7885
X1880 241 1 232 210 12 11 97 11 FA_X1 $T=1000 9400 1 0 $X=885 $Y=7885
X1881 128 2 52 241 12 11 98 11 FA_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X1882 69 164 211 132 12 11 242 11 FA_X1 $T=2330 9400 0 0 $X=2215 $Y=9285
X1883 70 135 186 242 12 11 189 11 FA_X1 $T=4040 12200 0 0 $X=3925 $Y=12085
X1884 211 165 243 187 12 11 99 11 FA_X1 $T=9360 9400 0 0 $X=9245 $Y=9285
X1885 244 3 84 253 12 11 100 11 FA_X1 $T=15820 9400 0 180 $X=12665 $Y=7885
X1886 129 142 189 143 12 11 102 11 FA_X1 $T=12780 12200 0 0 $X=12665 $Y=12085
X1887 130 168 188 244 12 11 101 11 FA_X1 $T=17150 9400 1 180 $X=13995 $Y=9285
X1888 164 166 213 246 12 11 264 11 FA_X1 $T=15060 12200 1 0 $X=14945 $Y=10685
X1889 188 167 212 254 12 11 245 11 FA_X1 $T=15820 9400 1 0 $X=15705 $Y=7885
X1890 19 169 234 245 12 11 103 11 FA_X1 $T=18860 9400 1 0 $X=18745 $Y=7885
X1891 168 214 233 255 12 11 234 11 FA_X1 $T=18860 9400 0 0 $X=18745 $Y=9285
X1892 186 85 54 264 12 11 104 11 FA_X1 $T=18860 12200 0 0 $X=18745 $Y=12085
X1893 119 86 72 145 12 11 169 11 FA_X1 $T=24560 12200 0 180 $X=21405 $Y=10685
X1894 118 190 235 215 12 11 105 11 FA_X1 $T=22280 9400 0 0 $X=22165 $Y=9285
X1895 120 191 192 216 12 11 106 11 FA_X1 $T=27980 12200 1 0 $X=27865 $Y=10685
X1896 26 87 217 218 12 11 107 11 FA_X1 $T=30070 9400 1 0 $X=29955 $Y=7885
X1897 56 136 55 133 12 11 25 11 FA_X1 $T=33300 12200 1 180 $X=30145 $Y=12085
X1898 218 236 137 134 12 11 57 11 FA_X1 $T=33110 9400 1 0 $X=32995 $Y=7885
X1899 217 170 193 247 12 11 194 11 FA_X1 $T=33870 12200 0 0 $X=33755 $Y=12085
X1900 73 171 195 88 12 11 74 11 FA_X1 $T=35200 9400 0 0 $X=35085 $Y=9285
X1901 171 172 256 196 12 11 5 11 FA_X1 $T=36150 9400 1 0 $X=36035 $Y=7885
X1902 131 6 58 194 12 11 108 11 FA_X1 $T=40520 12200 1 180 $X=37365 $Y=12085
X1903 172 173 248 237 12 11 197 11 FA_X1 $T=38810 9400 0 0 $X=38695 $Y=9285
X1904 195 89 138 198 12 11 109 11 FA_X1 $T=40520 12200 0 0 $X=40405 $Y=12085
X1905 198 262 219 257 12 11 249 11 FA_X1 $T=42230 12200 1 0 $X=42115 $Y=10685
X1906 121 90 249 197 12 11 32 11 FA_X1 $T=42800 9400 0 0 $X=42685 $Y=9285
X1907 122 174 91 259 12 11 36 11 FA_X1 $T=45270 12200 1 0 $X=45155 $Y=10685
X1908 38 175 199 258 12 11 40 11 FA_X1 $T=48500 9400 1 0 $X=48385 $Y=7885
X1909 123 223 144 201 12 11 110 11 FA_X1 $T=51920 9400 1 0 $X=51805 $Y=7885
X1910 259 176 200 51 12 11 201 11 FA_X1 $T=56670 12200 1 180 $X=53515 $Y=12085
X1911 174 7 220 221 12 11 111 11 FA_X1 $T=54390 12200 1 0 $X=54275 $Y=10685
X1912 220 139 203 202 12 11 76 11 FA_X1 $T=57240 12200 0 0 $X=57125 $Y=12085
X1913 221 177 222 204 12 11 77 11 FA_X1 $T=58950 9400 0 0 $X=58835 $Y=9285
X1914 124 43 225 92 12 11 41 11 FA_X1 $T=63510 12200 0 180 $X=60355 $Y=10685
X1915 179 178 224 226 12 11 112 11 FA_X1 $T=62370 9400 1 0 $X=62255 $Y=7885
X1916 223 179 250 140 12 11 225 11 FA_X1 $T=62370 9400 0 0 $X=62255 $Y=9285
X1917 250 180 227 260 12 11 113 11 FA_X1 $T=63510 12200 1 0 $X=63395 $Y=10685
X1918 224 141 93 94 12 11 251 11 FA_X1 $T=72250 12200 1 180 $X=69095 $Y=12085
X1919 125 95 182 251 12 11 114 11 FA_X1 $T=69400 9400 1 0 $X=69285 $Y=7885
X1920 178 181 252 183 12 11 182 11 FA_X1 $T=69590 9400 0 0 $X=69475 $Y=9285
X1921 64 205 238 261 12 11 115 11 FA_X1 $T=73010 9400 1 0 $X=72895 $Y=7885
X1922 116 228 206 207 12 11 229 11 FA_X1 $T=77000 12200 1 180 $X=73845 $Y=12085
X1923 48 184 230 208 12 11 239 11 FA_X1 $T=77000 12200 1 0 $X=76885 $Y=10685
X1924 79 8 239 229 12 11 185 11 FA_X1 $T=78140 9400 0 0 $X=78025 $Y=9285
.ENDS
***************************************
.SUBCKT ICV_24 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96
** N=284 EP=95 IP=3265 FDC=1916
M0 30 152 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=36675 $Y=1090 $D=1
M1 16 152 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=36865 $Y=1090 $D=1
M2 30 152 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37055 $Y=1090 $D=1
M3 16 152 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37245 $Y=1090 $D=1
M4 30 153 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37435 $Y=1090 $D=1
M5 16 153 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37625 $Y=1090 $D=1
M6 30 153 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=37815 $Y=1090 $D=1
M7 16 153 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=38005 $Y=1090 $D=1
M8 16 155 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=38425 $Y=1090 $D=1
M9 30 155 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38615 $Y=1090 $D=1
M10 16 155 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38805 $Y=1090 $D=1
M11 30 155 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=38995 $Y=1090 $D=1
M12 16 157 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39185 $Y=1090 $D=1
M13 30 157 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39375 $Y=1090 $D=1
M14 16 157 30 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=39565 $Y=1090 $D=1
M15 30 157 16 284 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=39755 $Y=1090 $D=1
M16 30 152 154 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=36675 $Y=1680 $D=0
M17 154 152 30 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=36865 $Y=1680 $D=0
M18 30 152 154 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37055 $Y=1680 $D=0
M19 154 152 30 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37245 $Y=1680 $D=0
M20 156 153 154 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37435 $Y=1680 $D=0
M21 154 153 156 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37625 $Y=1680 $D=0
M22 156 153 154 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=37815 $Y=1680 $D=0
M23 154 153 156 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=38005 $Y=1680 $D=0
M24 156 155 158 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=38425 $Y=1680 $D=0
M25 158 155 156 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38615 $Y=1680 $D=0
M26 156 155 158 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38805 $Y=1680 $D=0
M27 158 155 156 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=38995 $Y=1680 $D=0
M28 17 157 158 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39185 $Y=1680 $D=0
M29 158 157 17 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39375 $Y=1680 $D=0
M30 17 157 158 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=39565 $Y=1680 $D=0
M31 158 157 17 17 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=39755 $Y=1680 $D=0
X1595 177 110 16 17 152 284 AND2_X1 $T=30640 1000 0 0 $X=30525 $Y=885
X1596 196 125 16 17 234 284 AND2_X1 $T=55150 1000 0 0 $X=55035 $Y=885
X1597 214 143 16 17 162 284 AND2_X1 $T=79090 1000 0 0 $X=78975 $Y=885
X1711 160 121 230 117 16 17 OAI21_X1 $T=46980 3800 0 180 $X=46105 $Y=2285
X1712 208 139 270 136 16 17 OAI21_X1 $T=69210 3800 1 0 $X=69095 $Y=2285
X1779 183 16 17 181 16 INV_X1 $T=34630 3800 0 180 $X=34135 $Y=2285
X1780 186 16 17 262 284 INV_X1 $T=41090 1000 1 180 $X=40595 $Y=885
X1781 198 16 17 266 16 INV_X1 $T=60660 3800 0 180 $X=60165 $Y=2285
X1782 204 16 17 268 284 INV_X1 $T=66550 1000 1 180 $X=66055 $Y=885
X1783 219 16 17 220 16 INV_X1 $T=81560 3800 1 0 $X=81445 $Y=2285
X1894 110 175 279 16 17 227 16 HA_X1 $T=27980 3800 0 0 $X=27865 $Y=3685
X1895 68 227 226 16 17 28 16 HA_X1 $T=30070 6600 0 180 $X=28055 $Y=5085
X1896 151 182 112 16 17 175 16 HA_X1 $T=35010 3800 0 0 $X=34895 $Y=3685
X1897 159 191 252 16 17 182 16 HA_X1 $T=42230 3800 0 0 $X=42115 $Y=3685
X1898 160 192 283 16 17 191 16 HA_X1 $T=46030 3800 1 180 $X=44015 $Y=3685
X1899 125 254 126 16 17 192 16 HA_X1 $T=55720 3800 0 0 $X=55605 $Y=3685
X1900 240 202 132 16 17 254 16 HA_X1 $T=62370 3800 0 0 $X=62255 $Y=3685
X1901 134 203 137 16 17 132 16 HA_X1 $T=64840 3800 0 0 $X=64725 $Y=3685
X1902 208 212 140 16 17 137 16 HA_X1 $T=69970 3800 1 0 $X=69855 $Y=2285
X1903 143 34 142 16 17 140 284 HA_X1 $T=79090 1000 1 180 $X=77075 $Y=885
X1904 244 89 144 16 17 141 16 HA_X1 $T=80610 3800 1 180 $X=78595 $Y=3685
X1973 17 150 70 280 16 16 XOR2_X1 $T=33110 6600 1 0 $X=32995 $Y=5085
X1974 17 186 231 190 16 284 XOR2_X1 $T=43940 1000 1 180 $X=42685 $Y=885
X1975 17 120 232 230 16 16 XOR2_X1 $T=54010 3800 1 0 $X=53895 $Y=2285
X1976 17 238 236 239 16 16 XOR2_X1 $T=59330 3800 0 180 $X=58075 $Y=2285
X1977 17 204 209 269 16 16 XOR2_X1 $T=67500 3800 0 180 $X=66245 $Y=2285
X1978 17 138 210 270 16 284 XOR2_X1 $T=69400 1000 0 0 $X=69285 $Y=885
X1979 17 242 245 246 16 284 XOR2_X1 $T=83080 1000 0 0 $X=82965 $Y=885
X1982 151 16 180 183 17 284 NAND2_X1 $T=34820 1000 1 180 $X=34135 $Y=885
X1983 159 16 118 116 17 16 NAND2_X1 $T=40520 3800 0 180 $X=39835 $Y=2285
X1984 160 16 121 117 17 284 NAND2_X1 $T=45270 1000 0 0 $X=45155 $Y=885
X1985 240 16 129 198 17 16 NAND2_X1 $T=60090 3800 0 0 $X=59975 $Y=3685
X1986 134 16 135 133 17 16 NAND2_X1 $T=63320 3800 1 0 $X=63205 $Y=2285
X1987 208 16 139 136 17 284 NAND2_X1 $T=68830 1000 0 0 $X=68715 $Y=885
X1988 244 16 218 219 17 16 NAND2_X1 $T=82130 3800 1 180 $X=81445 $Y=3685
X1989 37 17 36 102 16 16 NOR2_X1 $T=2140 3800 0 0 $X=2025 $Y=3685
X1990 37 17 32 101 16 16 NOR2_X1 $T=2330 3800 1 0 $X=2215 $Y=2285
X1991 20 17 36 163 16 16 NOR2_X1 $T=5370 3800 1 0 $X=5255 $Y=2285
X1992 20 17 18 164 16 16 NOR2_X1 $T=5370 3800 0 0 $X=5255 $Y=3685
X1993 19 17 18 221 16 284 NOR2_X1 $T=6890 1000 1 180 $X=6205 $Y=885
X1994 19 17 25 222 16 16 NOR2_X1 $T=6890 6600 0 180 $X=6205 $Y=5085
X1995 20 17 32 165 16 16 NOR2_X1 $T=8220 3800 1 0 $X=8105 $Y=2285
X1996 37 17 21 103 16 16 NOR2_X1 $T=8410 3800 0 0 $X=8295 $Y=3685
X1997 38 17 25 47 16 16 NOR2_X1 $T=11450 6600 0 0 $X=11335 $Y=6485
X1998 19 17 36 166 16 284 NOR2_X1 $T=12400 1000 1 180 $X=11715 $Y=885
X1999 38 17 18 104 16 16 NOR2_X1 $T=12020 6600 1 0 $X=11905 $Y=5085
X2000 31 17 23 24 16 16 NOR2_X1 $T=12020 6600 0 0 $X=11905 $Y=6485
X2001 31 17 25 147 16 16 NOR2_X1 $T=12590 6600 1 0 $X=12475 $Y=5085
X2002 40 17 23 273 16 16 NOR2_X1 $T=14680 6600 1 180 $X=13995 $Y=6485
X2003 110 17 177 179 16 16 NOR2_X1 $T=31210 3800 0 180 $X=30525 $Y=2285
X2004 152 17 179 178 16 284 NOR2_X1 $T=31400 1000 0 0 $X=31285 $Y=885
X2005 31 17 18 29 16 16 NOR2_X1 $T=33110 6600 0 0 $X=32995 $Y=6485
X2006 151 17 180 113 16 284 NOR2_X1 $T=33680 1000 0 0 $X=33565 $Y=885
X2007 181 17 113 280 16 16 NOR2_X1 $T=34250 3800 0 180 $X=33565 $Y=2285
X2008 40 17 25 42 16 16 NOR2_X1 $T=35200 6600 0 0 $X=35085 $Y=6485
X2009 183 17 179 153 16 284 NOR2_X1 $T=35960 1000 0 0 $X=35845 $Y=885
X2010 159 17 118 114 16 16 NOR2_X1 $T=39950 3800 0 0 $X=39835 $Y=3685
X2011 160 17 121 188 16 284 NOR2_X1 $T=45270 1000 1 180 $X=44585 $Y=885
X2012 38 17 21 123 16 16 NOR2_X1 $T=51160 6600 0 180 $X=50475 $Y=5085
X2013 40 17 36 194 16 16 NOR2_X1 $T=53060 6600 1 180 $X=52375 $Y=6485
X2014 31 17 32 282 16 16 NOR2_X1 $T=54390 6600 1 0 $X=54275 $Y=5085
X2015 125 17 196 195 16 284 NOR2_X1 $T=54580 1000 0 0 $X=54465 $Y=885
X2016 234 17 195 237 16 16 NOR2_X1 $T=57620 3800 1 0 $X=57505 $Y=2285
X2017 266 17 130 239 16 284 NOR2_X1 $T=60280 1000 1 180 $X=59595 $Y=885
X2018 240 17 129 130 16 16 NOR2_X1 $T=60660 3800 0 0 $X=60545 $Y=3685
X2019 198 17 195 199 16 16 NOR2_X1 $T=61420 3800 1 0 $X=61305 $Y=2285
X2020 134 17 135 131 16 16 NOR2_X1 $T=64840 3800 1 180 $X=64155 $Y=3685
X2021 208 17 139 206 16 16 NOR2_X1 $T=69210 3800 0 180 $X=68525 $Y=2285
X2022 44 17 21 271 16 16 NOR2_X1 $T=69780 6600 0 0 $X=69665 $Y=6485
X2023 143 17 214 145 16 16 NOR2_X1 $T=79280 3800 0 180 $X=78595 $Y=2285
X2024 162 17 145 215 16 16 NOR2_X1 $T=80040 3800 1 0 $X=79925 $Y=2285
X2025 219 17 145 216 16 16 NOR2_X1 $T=80610 6600 1 0 $X=80495 $Y=5085
X2026 244 17 218 146 16 16 NOR2_X1 $T=83080 3800 0 0 $X=82965 $Y=3685
X2027 220 17 146 246 16 284 NOR2_X1 $T=84220 1000 0 0 $X=84105 $Y=885
X2028 262 116 150 114 16 17 16 AOI21_X1 $T=39950 3800 0 180 $X=39075 $Y=2285
X2029 116 117 155 187 16 17 284 AOI21_X1 $T=39950 1000 0 0 $X=39835 $Y=885
X2030 159 118 190 114 16 17 16 AOI21_X1 $T=41850 3800 0 180 $X=40975 $Y=2285
X2031 117 120 186 188 16 17 16 AOI21_X1 $T=42990 3800 1 0 $X=42875 $Y=2285
X2032 268 133 238 131 16 17 284 AOI21_X1 $T=63320 1000 0 0 $X=63205 $Y=885
X2033 134 135 269 131 16 17 16 AOI21_X1 $T=63890 3800 1 0 $X=63775 $Y=2285
X2034 133 136 200 205 16 17 284 AOI21_X1 $T=64080 1000 0 0 $X=63965 $Y=885
X2035 136 138 204 206 16 17 284 AOI21_X1 $T=68070 1000 1 180 $X=67195 $Y=885
X2036 74 13 242 15 16 17 16 AOI21_X1 $T=83080 6600 1 180 $X=82205 $Y=6485
X2037 13 14 217 51 16 17 16 AOI21_X1 $T=83080 6600 1 0 $X=82965 $Y=5085
X2038 120 17 188 187 16 157 284 NOR3_X1 $T=41850 1000 1 180 $X=40975 $Y=885
X2039 138 17 206 205 16 241 284 NOR3_X1 $T=67310 1000 1 180 $X=66435 $Y=885
X2040 16 178 69 111 17 16 XNOR2_X1 $T=31590 3800 1 0 $X=31475 $Y=2285
X2041 16 237 235 127 17 284 XNOR2_X1 $T=58000 1000 1 180 $X=56745 $Y=885
X2042 16 215 211 243 17 284 XNOR2_X1 $T=79850 1000 0 0 $X=79735 $Y=885
X2043 179 113 114 16 17 187 OR3_X1 $T=36720 3800 1 0 $X=36605 $Y=2285
X2044 195 130 131 16 17 205 OR3_X1 $T=62370 3800 1 0 $X=62255 $Y=2285
X2045 145 146 15 16 17 51 OR3_X1 $T=83840 6600 1 0 $X=83725 $Y=5085
X2046 150 181 16 111 180 151 17 OAI22_X1 $T=32730 3800 1 0 $X=32615 $Y=2285
X2047 238 266 16 127 129 240 17 OAI22_X1 $T=59330 3800 1 0 $X=59215 $Y=2285
X2048 242 220 16 243 218 244 17 OAI22_X1 $T=82320 3800 1 0 $X=82205 $Y=2285
X2050 236 17 235 232 231 50 16 16 NOR4_X1 $T=56100 3800 0 180 $X=55035 $Y=2285
X2051 241 17 200 199 234 120 16 284 NOR4_X1 $T=61990 1000 1 180 $X=60925 $Y=885
X2052 245 17 211 210 209 45 16 284 NOR4_X1 $T=73580 1000 1 180 $X=72515 $Y=885
X2053 46 17 217 216 162 138 16 16 NOR4_X1 $T=81560 3800 1 180 $X=80495 $Y=3685
X2054 71 101 163 221 17 16 248 284 FA_X1 $T=1000 1000 0 0 $X=885 $Y=885
X2055 67 102 164 222 17 16 258 16 FA_X1 $T=2330 6600 1 0 $X=2215 $Y=5085
X2056 72 52 258 75 17 16 259 16 FA_X1 $T=8410 6600 0 0 $X=8295 $Y=6485
X2057 247 103 165 166 17 16 223 284 FA_X1 $T=11830 1000 1 180 $X=8675 $Y=885
X2058 105 278 247 90 17 16 106 16 FA_X1 $T=12020 6600 0 180 $X=8865 $Y=5085
X2059 278 104 147 273 17 16 249 16 FA_X1 $T=12780 3800 0 0 $X=12665 $Y=3685
X2060 39 169 167 259 17 16 108 284 FA_X1 $T=13540 1000 0 0 $X=13425 $Y=885
X2061 73 224 54 96 17 16 167 16 FA_X1 $T=14870 6600 1 0 $X=14755 $Y=5085
X2062 224 53 248 55 17 16 225 16 FA_X1 $T=15820 3800 0 0 $X=15705 $Y=3685
X2063 168 26 249 223 17 16 109 284 FA_X1 $T=16580 1000 0 0 $X=16465 $Y=885
X2064 27 105 171 76 17 16 260 16 FA_X1 $T=17910 6600 1 0 $X=17795 $Y=5085
X2065 48 1 170 260 17 16 148 16 FA_X1 $T=18860 3800 0 0 $X=18745 $Y=3685
X2066 169 56 250 168 17 16 176 284 FA_X1 $T=19620 1000 0 0 $X=19505 $Y=885
X2067 170 106 174 77 17 16 107 16 FA_X1 $T=20950 6600 1 0 $X=20835 $Y=5085
X2068 251 107 172 225 17 16 173 16 FA_X1 $T=22280 3800 0 0 $X=22165 $Y=3685
X2069 171 84 41 57 17 16 174 16 FA_X1 $T=22280 6600 0 0 $X=22165 $Y=6485
X2070 226 108 251 148 17 16 177 284 FA_X1 $T=22660 1000 0 0 $X=22545 $Y=885
X2071 279 173 176 149 17 16 180 284 FA_X1 $T=27600 1000 0 0 $X=27485 $Y=885
X2072 149 109 228 189 17 16 115 16 FA_X1 $T=30070 6600 1 0 $X=29955 $Y=5085
X2073 250 2 92 91 17 16 228 16 FA_X1 $T=30070 6600 0 0 $X=29955 $Y=6485
X2074 172 58 184 78 17 16 261 16 FA_X1 $T=35770 6600 0 0 $X=35655 $Y=6485
X2075 112 115 185 261 17 16 118 16 FA_X1 $T=36910 3800 0 0 $X=36795 $Y=3685
X2076 184 3 59 229 17 16 119 16 FA_X1 $T=38810 6600 0 0 $X=38695 $Y=6485
X2077 185 119 49 281 17 16 283 16 FA_X1 $T=42230 6600 1 0 $X=42115 $Y=5085
X2078 189 60 85 61 17 16 263 16 FA_X1 $T=42230 6600 0 0 $X=42115 $Y=6485
X2079 229 4 253 79 17 16 161 16 FA_X1 $T=45270 6600 0 0 $X=45155 $Y=6485
X2080 252 122 193 263 17 16 121 284 FA_X1 $T=48880 1000 1 180 $X=45725 $Y=885
X2081 281 161 93 80 17 16 264 16 FA_X1 $T=46030 3800 0 0 $X=45915 $Y=3685
X2082 253 123 282 194 17 16 265 16 FA_X1 $T=48310 6600 0 0 $X=48195 $Y=6485
X2083 193 5 62 274 17 16 124 16 FA_X1 $T=50970 3800 1 0 $X=50855 $Y=2285
X2084 122 124 264 275 17 16 196 284 FA_X1 $T=51540 1000 0 0 $X=51425 $Y=885
X2085 274 6 265 63 17 16 233 16 FA_X1 $T=52680 3800 0 0 $X=52565 $Y=3685
X2086 275 7 197 94 17 16 128 16 FA_X1 $T=55910 6600 0 0 $X=55795 $Y=6485
X2087 126 128 233 81 17 16 129 16 FA_X1 $T=57050 6600 1 0 $X=56935 $Y=5085
X2088 197 8 43 17 17 16 201 16 FA_X1 $T=58950 6600 0 0 $X=58835 $Y=6485
X2089 202 9 201 267 17 16 135 16 FA_X1 $T=62370 6600 0 0 $X=62255 $Y=6485
X2090 267 10 255 86 17 16 207 16 FA_X1 $T=65410 6600 0 0 $X=65295 $Y=6485
X2091 203 207 33 95 17 16 139 16 FA_X1 $T=66740 3800 0 0 $X=66625 $Y=3685
X2092 255 276 277 82 17 16 257 16 FA_X1 $T=69780 3800 0 0 $X=69665 $Y=3685
X2093 276 64 271 87 17 16 256 16 FA_X1 $T=72820 6600 0 0 $X=72705 $Y=6485
X2094 212 141 272 257 17 16 214 16 FA_X1 $T=75670 3800 1 0 $X=75555 $Y=2285
X2095 272 256 35 65 17 16 144 16 FA_X1 $T=75670 3800 0 0 $X=75555 $Y=3685
X2096 277 11 88 83 17 16 213 16 FA_X1 $T=75860 6600 0 0 $X=75745 $Y=6485
X2097 142 12 213 66 17 16 218 16 FA_X1 $T=78900 6600 0 0 $X=78785 $Y=6485
.ENDS
***************************************
.SUBCKT FloatingPointMultiplierSingle VSS VDD result[31] result[30] result[29] result[27] result[26] result[23] result[25] result[22] result[24] result[21] result[20] inputA[16] inputB[16] result[19] inputB[13] result[18] inputB[11] inputB[9]
+ inputB[14] inputA[14] inputA[8] result[17] inputA[11] inputA[6] inputA[10] inputA[12] inputA[9] inputA[7] inputA[13] result[16] result[15] result[14] result[13] result[12] en reset result[11] clk
+ result[0] inputB[31] inputB[17] inputB[25] inputB[28] inputA[20] inputB[18] inputB[3] inputA[1] inputA[2] inputA[3] inputA[0] result[28] result[10] result[6] result[7] result[9] OF result[4] result[2]
+ result[1] result[8] inputB[22] inputB[29] inputB[26] inputB[23] result[5] result[3] inputA[25] inputA[17] inputA[30] inputA[27] inputA[21] inputB[21] inputB[15] inputA[29] inputA[26] inputA[28] inputA[22] inputB[20]
+ inputA[24] inputA[23] inputA[31] inputB[27] inputB[24] inputB[19] inputB[30] inputB[4] inputA[4] inputB[5] inputB[6] inputA[5] inputB[8] inputA[15] inputB[7] inputA[18] inputB[10] inputA[19] inputB[12] inputB[2]
+ inputB[1] inputB[0]
** N=881 EP=102 IP=2108 FDC=22878
X0 86 11 16 19 20 27 35 36 inputB[16] inputA[16] 40 10 44 inputB[11] inputB[14] inputB[9] 53 inputA[14] 56 inputA[13]
+ inputA[12] inputA[11] inputA[10] inputA[9] inputA[8] 68 71 72 74 77 reset clk 7 VDD VSS result[30] result[29] result[26] result[22] 39
+ 47 result[18] 70 inputA[7] 69 79 result[13] 835 13 28 30 37 41 result[19] 6 91 93 78 85 result[11]
+ en result[9] result[28] result[24] 34 50 63 66 92 result[15] result[10] result[31] 31 result[20] 60 9 result[27] result[23] result[25] result[21]
+ result[17] result[16] result[14] result[12] 22 14 18 25 33 81 83 76 32
+ ICV_10 $T=0 0 0 0 $X=0 $Y=79285
X1 68 16 101 106 110 149 35 113 119 120 53 125 inputB[13] 131 134 135 139 69 inputA[6] 161
+ 175 152 156 158 160 155 162 166 168 167 169 86 VDD VSS 99 13 31 7 129 836
+ 145 147 157 30 10 148 9 835 18 25 118 114 116 117 124 122 34 862 128 871
+ 56 137 151 76 78 164 83 172 result[8] result[0] result[6] 105 115 126 44 127 94 70 153 150
+ 102 123 37 130 142 11 14 19 20 27 36 870 132 873 71 72 154 74 77 163
+ 79 81 170 173 171 96 95 136 144 143 146 result[7] 856 39 41 47 50 63 60 66
+ 85 22 32 133 138 100 103 111 112 28 121 33 97 98 104 107 109 108 140 141
+ 159 165 40
+ ICV_11 $T=0 0 0 0 $X=0 $Y=73685
X2 inputA[31] inputB[31] 53 96 874 180 182 98 101 181 183 106 109 105 107 110 108 252 185 186
+ 189 190 199 132 131 137 207 149 214 148 227 223 158 160 162 320 233 234 236 167
+ 241 838 170 86 7 VSS 99 104 184 864 VDD 111 30 187 188 124 119 120 192 125
+ 128 127 133 204 135 139 652 577 150 220 165 243 10 244 result[4] 35 70 861 179 114
+ 112 115 193 122 191 194 197 129 201 136 863 290 155 222 225 865 230 240 238 result[2]
+ OF 16 113 117 121 123 116 198 134 138 210 157 156 235 237 239 result[3] result[1] 206 208
+ 245 211 212 242 218 154 856 97 102 141 140 147 153 175 159 231 213 169 177 173
+ 171 100 103 13 126 130 142 145 151 152 164 876 166 118 200 203 209 221 875 202
+ 215 224 226 163 232 168 837 216 217 195 196 205 219 228 229
+ ICV_12 $T=0 0 0 0 $X=0 $Y=68085
X3 inputB[29] 53 inputB[23] inputB[26] inputB[22] inputB[25] inputB[17] 68 261 264 839 281 91 144 308 300 314 840 172 86
+ 2 7 VDD VSS 182 181 254 192 190 265 273 278 279 6 283 286 288 287 305 284
+ 94 291 143 215 330 219 226 316 233 336 239 337 216 257 285 280 205 211 92 146
+ 298 322 309 93 222 310 229 301 312 328 183 259 188 189 262 877 837 212 313 793
+ 227 388 236 329 867 235 241 878 258 866 260 268 269 272 274 277 276 296 293 294
+ 319 323 324 327 334 177 253 110 191 195 193 196 198 200 199 202 204 208 210 295
+ 224 232 230 325 234 238 243 838 292 297 306 794 311 318 result[5] 248 249 251 194 179
+ 109 106 255 108 113 187 197 203 206 209 218 228 223 240 256 275 289 299 304 307
+ 321 231 857 332 247 263 266 267 271 282 303 315 333 302 326 335 317 237 331 270
+ ICV_13 $T=0 0 0 0 $X=0 $Y=62485
X4 inputA[29] inputA[30] inputB[27] inputB[21] inputA[28] inputB[30] 68 inputA[17] inputB[28] inputB[24] inputB[15] 53 inputA[25] inputA[26] inputB[20] inputA[24] inputA[23] inputA[22] inputA[21] inputB[19]
+ 350 345 264 304 368 VDD 841 339 386 373 395 401 VSS 207 2 7 70 341 248 180
+ 255 107 347 348 349 256 351 357 278 353 284 355 312 367 265 359 266 364 370 269
+ 201 378 346 362 272 273 369 277 286 863 873 299 399 301 217 380 308 865 94 221
+ 381 315 358 285 379 321 326 338 394 390 404 305 406 337 inputA[27] 253 98 101 184 257
+ 259 262 263 267 839 365 275 276 281 282 288 374 245 293 213 303 220 387 314 398
+ 875 298 328 331 878 861 352 189 260 185 344 356 95 862 280 871 274 295 287 400
+ 385 313 319 318 405 333 334 354 360 283 292 306 794 311 391 392 325 396 397 402
+ 484 407 249 343 874 186 258 261 268 271 279 294 844 289 291 252 296 307 382 383
+ 793 225 324 323 332 336 361 377 384 389 836 254 251 270 290 162 302 317 327 857
+ 244 366 6 363 376 393 408 403 372 309 375 858 371 297 316
+ ICV_16 $T=0 0 0 0 $X=0 $Y=51285
X5 inputB[3] inputB[4] inputB[6] inputA[20] inputA[18] inputB[18] inputA[19] inputA[15] inputB[7] 53 68 inputB[10] inputB[8] inputA[5] inputB[12] 349 358 301 412 828
+ 567 872 437 413 876 304 475 424 VDD 247 VSS 70 344 7 322 364 414 285 421 420
+ 373 416 422 357 308 426 415 284 278 398 431 312 399 363 365 434 419 338 378 447
+ 380 452 453 329 175 382 320 330 391 405 384 472 310 471 393 369 379 381 469 346
+ 479 396 406 362 inputB[5] 351 367 425 423 354 313 361 842 148 829 442 370 446 376 242
+ 458 160 383 462 387 476 298 843 840 407 880 397 355 360 348 305 350 352 866 877
+ 868 158 867 459 482 464 394 467 392 480 395 356 214 436 445 448 454 457 879 389
+ 477 404 353 427 429 359 366 841 371 374 449 300 461 466 470 390 486 408 403 859
+ 418 432 433 489 440 443 463 478 484 341 411 343 870 441 347 345 368 372 161 375
+ 386 388 401 335 417 465 474 487 864 430 438 450 377 456 460 488 468 385 473 483
+ 485 428 409 455 402 451 435 439 444 481
+ ICV_17 $T=0 0 0 0 $X=0 $Y=40085
X6 inputB[1] inputB[0] 53 inputA[4] 512 509 68 524 527 557 461 469 511 549 550 551 556 339 VSS VDD
+ 7 338 373 285 417 364 415 416 308 419 322 424 313 346 422 423 398 379 384 431
+ 380 399 310 378 381 420 529 437 414 520 438 842 530 443 449 444 454 452 533 534
+ 536 456 539 459 304 543 465 515 362 370 278 312 301 476 479 369 298 475 477 367
+ 554 482 487 558 486 400 inputB[2] 70 330 436 522 442 446 590 531 305 521 468 485 555
+ 411 412 494 497 498 502 503 501 435 504 507 508 433 441 532 440 513 537 462 491
+ 495 421 425 357 516 528 829 540 466 470 472 548 478 480 492 493 428 510 448 445
+ 453 451 455 545 546 458 473 474 843 488 483 833 538 535 413 430 450 447 457 460
+ 471 880 427 506 429 525 464 490 418 500 426 432 517 518 519 523 526 542 467 544
+ 553 496 499 541 845 547 552 505 439 463
+ ICV_18 $T=0 0 0 0 $X=0 $Y=30180
X7 846 504 580 278 527 587 540 597 602 833 VSS VDD 338 491 373 422 367 416 308 506
+ 500 502 384 511 507 574 515 572 514 419 517 312 284 526 378 513 529 534 521 535
+ 592 591 400 844 595 414 380 544 547 304 298 606 301 481 285 379 558 305 495 330
+ 424 369 362 523 582 588 541 542 346 420 364 598 548 549 370 550 610 551 554 561
+ 415 563 310 399 569 570 575 576 581 583 599 600 543 845 858 417 611 879 494 498
+ 579 586 537 546 559 564 565 496 409 571 573 512 520 539 524 605 552 555 585 596
+ 601 594 556 497 505 509 584 536 528 553 560 493 510 525 603 589 538 848 849 322
+ 398 847 492 503 566 562 508 593 604 609 568 578 608 501 545 607
+ ICV_19 $T=0 0 0 0 $X=0 $Y=24685
X8 569 513 571 636 581 68 601 606 651 610 4 VSS VDD 338 373 285 415 562 298 566
+ 398 511 378 574 369 515 570 850 434 577 310 399 522 525 584 362 313 304 301 521
+ 308 379 594 593 469 370 648 322 849 607 417 572 613 420 560 414 626 499 384 568
+ 575 516 634 489 631 330 582 586 588 589 557 284 848 531 597 602 604 380 609 381
+ 305 608 846 622 628 632 633 624 635 214 868 519 532 643 598 647 653 654 416 851
+ 559 616 564 623 621 619 637 638 640 644 605 656 490 614 618 620 578 518 580 579
+ 530 587 590 603 658 657 630 655 834 639 567 533 659 629 561 617 563 625 854 583
+ 649 615 585 642 592 596 646 650 627 576 573 645 599 600 612 565 641 611
+ ICV_20 $T=0 0 0 0 $X=0 $Y=19085
X9 663 667 381 570 872 inputA[1] 68 inputA[2] inputA[3] 398 417 420 656 710 4 VSS VDD 416 298 419
+ 330 313 628 625 627 369 574 362 572 676 678 634 636 310 424 399 70 308 521 469
+ 380 690 384 322 285 591 513 422 595 511 414 699 700 515 651 704 653 705 inputA[0] 620
+ 379 378 633 677 685 642 305 540 694 644 415 703 650 652 707 657 712 658 626 674
+ 675 679 635 638 687 640 643 692 693 755 645 646 698 647 648 649 701 711 881 706
+ 869 853 834 708 852 614 664 695 696 655 851 662 621 616 617 666 671 670 680 682
+ 639 683 641 691 697 702 673 850 681 686 709 689 847 615 619 629 631 632 637 661
+ 654 659 618 665 668 669 688 622 630 672
+ ICV_22 $T=0 0 0 0 $X=0 $Y=13485
X10 714 662 722 469 744 683 694 705 706 712 VSS VDD 285 415 330 313 424 726 399 310
+ 380 419 398 734 735 513 384 298 417 322 749 511 688 379 751 414 748 521 752 758
+ 416 698 570 572 515 422 769 771 710 692 613 373 671 678 730 739 682 308 695 696
+ 574 766 764 768 855 775 708 612 852 718 673 733 741 750 759 760 420 772 773 853
+ 860 777 721 670 672 680 681 685 687 690 697 702 703 704 709 716 663 719 720 725
+ 667 728 727 724 736 737 743 747 754 757 761 762 765 774 767 869 729 732 731 745
+ 746 753 756 763 770 776 661 623 669 742 715 679 740 717 675 738 686 693 699 701
+ 723 666 691 674
+ ICV_23 $T=0 0 0 0 $X=0 $Y=7885
X11 727 737 739 748 749 752 756 759 758 761 768 773 855 853 775 VSS VDD 414 298 308
+ 415 422 721 416 724 668 676 738 872 330 417 700 765 707 420 305 322 665 313 731
+ 740 760 384 881 860 722 723 743 711 777 719 720 726 735 728 729 741 744 745 746
+ 753 755 767 769 774 715 677 624 854 714 717 664 776 716 732 733 742 750 689 754
+ 764 771 730 747 762 766 770 772 718 736 734 751 757 763 725
+ ICV_24 $T=0 0 0 0 $X=0 $Y=0
.ENDS
***************************************
