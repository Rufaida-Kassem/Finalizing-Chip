* SPICE NETLIST
***************************************

*.CALIBRE ABORT_INFO SUPPLY_ERROR
.SUBCKT MGC_via1_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_1
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X2
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_AUTO_NDR_MGC_CLK_NDR_1.0w2.0s_via2_single_MA_north
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X4
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT CLKBUF_X3 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=8
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.0475e-14 PD=6.7e-07 PS=6e-07 $X=145 $Y=90 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=335 $Y=90 $D=1
M2 VSS 7 Z 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=525 $Y=90 $D=1
M3 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=715 $Y=90 $D=1
M4 VDD A 7 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 VDD 7 Z 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_3
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT FILLCELL_X8
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_4
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT DFF_X1 D CK VSS VDD Q 6 7
** N=22 EP=7 IP=0 FDC=28
M0 VSS 11 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=160 $Y=180 $D=1
M1 19 10 VSS 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.1e-14 PD=4.6e-07 PS=7e-07 $X=350 $Y=300 $D=1
M2 9 8 19 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.6e-14 AS=1.26e-14 PD=8.4e-07 PS=4.6e-07 $X=540 $Y=300 $D=1
M3 20 11 9 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=2.6e-14 PD=8.3e-07 PS=8.4e-07 $X=735 $Y=180 $D=1
M4 VSS D 20 6 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.395e-14 AS=3.85e-14 PD=8.3e-07 PS=8.3e-07 $X=925 $Y=180 $D=1
M5 10 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=3.395e-14 PD=6.3e-07 PS=8.3e-07 $X=1115 $Y=180 $D=1
M6 VSS CK 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1530 $Y=255 $D=1
M7 21 9 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1720 $Y=255 $D=1
M8 12 8 21 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.1e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1910 $Y=255 $D=1
M9 22 11 12 6 NMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.1e-14 PD=4.7e-07 PS=7e-07 $X=2100 $Y=300 $D=1
M10 VSS 14 22 6 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.305e-14 PD=7e-07 PS=4.7e-07 $X=2295 $Y=300 $D=1
M11 14 12 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=2485 $Y=255 $D=1
M12 VSS 12 QN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=2825 $Y=90 $D=1
M13 Q 14 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=3015 $Y=90 $D=1
M14 VDD 11 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=160 $Y=785 $D=0
M15 15 10 VDD 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.835e-14 PD=4.6e-07 PS=9.1e-07 $X=350 $Y=1010 $D=0
M16 9 11 15 7 PMOS_VTL L=5e-08 W=9e-08 AD=3.615e-14 AS=1.26e-14 PD=1.13e-06 PS=4.6e-07 $X=540 $Y=1010 $D=0
M17 16 8 9 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=3.615e-14 PD=1.12e-06 PS=1.13e-06 $X=735 $Y=765 $D=0
M18 VDD D 16 7 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.145e-14 AS=5.88e-14 PD=1.12e-06 PS=1.12e-06 $X=925 $Y=765 $D=0
M19 10 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.67e-14 AS=5.145e-14 PD=9.9e-07 PS=1.12e-06 $X=1115 $Y=870 $D=0
M20 VDD CK 11 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1530 $Y=870 $D=0
M21 17 9 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1720 $Y=870 $D=0
M22 12 11 17 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=2.835e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1910 $Y=870 $D=0
M23 18 8 12 7 PMOS_VTL L=5e-08 W=9e-08 AD=1.305e-14 AS=2.835e-14 PD=4.7e-07 PS=9.1e-07 $X=2100 $Y=1095 $D=0
M24 VDD 14 18 7 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.305e-14 PD=9.1e-07 PS=4.7e-07 $X=2295 $Y=1095 $D=0
M25 14 12 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=2485 $Y=870 $D=0
M26 VDD 12 QN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=2825 $Y=680 $D=0
M27 Q 14 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=3015 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=1 EP=0 IP=2 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKBUF_X1 A VSS VDD Z 5 6
** N=7 EP=6 IP=0 FDC=4
M0 VSS A 7 5 NMOS_VTL L=5e-08 W=9.5e-08 AD=2.03e-14 AS=9.975e-15 PD=6.7e-07 PS=4e-07 $X=165 $Y=160 $D=1
M1 Z 7 VSS 5 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.03e-14 PD=6e-07 PS=6.7e-07 $X=355 $Y=160 $D=1
M2 VDD A 7 6 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=3.3075e-14 PD=1.54e-06 PS=8.4e-07 $X=165 $Y=995 $D=0
M3 Z 7 VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=355 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via2_5
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT OR2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 8 A1 VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A1 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 9 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X32
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_HH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT AND2_X1 A1 A2 VSS VDD ZN 6 7
** N=9 EP=7 IP=0 FDC=6
M0 9 A1 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 9 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 ZN 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 8 A1 VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M4 VDD A2 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M5 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FILLCELL_X16
** N=4 EP=0 IP=0 FDC=0
*.CALIBRE ISOLATED NETS: VSS VDD
.ENDS
***************************************
.SUBCKT OAI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN B2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 9 B1 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=360 $Y=90 $D=1
M2 VSS A 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=550 $Y=90 $D=1
M3 10 B2 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M4 ZN B1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=360 $Y=680 $D=0
M5 VDD A ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=550 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT INV_X1 A VSS VDD ZN 5 6
** N=6 EP=6 IP=0 FDC=2
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.3575e-14 PD=1.04e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT HA_X1 S B A VSS VDD CO 7 8
** N=14 EP=8 IP=0 FDC=16
M0 13 B VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 S A 13 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS 10 S 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.48e-14 AS=5.81e-14 PD=1.12e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 10 B VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.48e-14 PD=7e-07 PS=1.12e-06 $X=760 $Y=90 $D=1
M4 VSS A 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=950 $Y=90 $D=1
M5 14 A 11 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1320 $Y=90 $D=1
M6 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=1510 $Y=90 $D=1
M7 CO 11 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1700 $Y=90 $D=1
M8 S B 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M9 9 A S 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M10 VDD 10 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.7725e-14 AS=8.82e-14 PD=1.55e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
M11 12 B VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.7725e-14 PD=9.1e-07 PS=1.55e-06 $X=760 $Y=870 $D=0
M12 10 A 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=950 $Y=870 $D=0
M13 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1320 $Y=870 $D=0
M14 VDD B 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=1510 $Y=870 $D=0
M15 CO 11 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1700 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT CLKGATETST_X1 SE E CK VDD VSS GCK 7 8
** N=20 EP=8 IP=0 FDC=24
M0 9 SE VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=205 $D=1
M1 VSS E 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.94e-14 PD=8.3e-07 PS=7e-07 $X=335 $Y=205 $D=1
M2 18 9 VSS 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=525 $Y=140 $D=1
M3 10 13 18 7 NMOS_VTL L=5e-08 W=2.75e-07 AD=2.915e-14 AS=3.85e-14 PD=9.1e-07 PS=8.3e-07 $X=715 $Y=140 $D=1
M4 19 11 10 7 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=2.915e-14 PD=4.6e-07 PS=9.1e-07 $X=945 $Y=300 $D=1
M5 VSS 12 19 7 NMOS_VTL L=5e-08 W=9e-08 AD=2.1e-14 AS=1.26e-14 PD=7e-07 PS=4.6e-07 $X=1135 $Y=300 $D=1
M6 11 13 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.1e-14 PD=6.3e-07 PS=7e-07 $X=1325 $Y=180 $D=1
M7 VSS 10 12 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1665 $Y=315 $D=1
M8 13 CK VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1855 $Y=315 $D=1
M9 20 CK 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=2240 $Y=295 $D=1
M10 VSS 10 20 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.835e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2430 $Y=295 $D=1
M11 GCK 14 VSS 7 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.835e-14 PD=6e-07 PS=7e-07 $X=2620 $Y=310 $D=1
M12 15 SE 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=890 $D=0
M13 VDD E 15 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=4.41e-14 PD=1.12e-06 PS=9.1e-07 $X=335 $Y=890 $D=0
M14 16 9 VDD 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=525 $Y=890 $D=0
M15 10 11 16 8 PMOS_VTL L=5e-08 W=4.2e-07 AD=3.93e-14 AS=5.88e-14 PD=1.2e-06 PS=1.12e-06 $X=715 $Y=890 $D=0
M16 17 13 10 8 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.93e-14 PD=4.6e-07 PS=1.2e-06 $X=945 $Y=990 $D=0
M17 VDD 12 17 8 PMOS_VTL L=5e-08 W=9e-08 AD=2.835e-14 AS=1.26e-14 PD=9.1e-07 PS=4.6e-07 $X=1135 $Y=990 $D=0
M18 11 13 VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=2.835e-14 PD=8.4e-07 PS=9.1e-07 $X=1325 $Y=990 $D=0
M19 VDD 10 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1665 $Y=870 $D=0
M20 13 CK VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1855 $Y=870 $D=0
M21 14 CK VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=2240 $Y=870 $D=0
M22 VDD 10 14 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2430 $Y=870 $D=0
M23 GCK 14 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2620 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT via1_7
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 98
** N=214 EP=91 IP=2606 FDC=1460
M0 124 37 37 211 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=77360 $Y=82290 $D=1
M1 37 125 124 211 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=77550 $Y=82290 $D=1
M2 37 128 126 211 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.395e-14 AS=2.205e-14 PD=8.3e-07 PS=6.3e-07 $X=77890 $Y=82290 $D=1
M3 205 124 37 211 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.85e-14 AS=3.395e-14 PD=8.3e-07 PS=8.3e-07 $X=78080 $Y=82290 $D=1
M4 129 128 205 211 NMOS_VTL L=5e-08 W=2.75e-07 AD=3.0125e-14 AS=3.85e-14 PD=8.7e-07 PS=8.3e-07 $X=78270 $Y=82290 $D=1
M5 206 126 129 211 NMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=3.0125e-14 PD=4.6e-07 PS=8.7e-07 $X=78480 $Y=82360 $D=1
M6 37 127 206 211 NMOS_VTL L=5e-08 W=9e-08 AD=3.58e-14 AS=1.26e-14 PD=1.12e-06 PS=4.6e-07 $X=78670 $Y=82360 $D=1
M7 127 129 37 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=3.58e-14 PD=1.11e-06 PS=1.12e-06 $X=78865 $Y=82290 $D=1
M8 37 129 127 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=79055 $Y=82290 $D=1
M9 37 131 128 211 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.69e-14 AS=3.36e-14 PD=1.14e-06 PS=7.4e-07 $X=79450 $Y=82290 $D=1
M10 207 131 37 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.69e-14 PD=1.11e-06 PS=1.14e-06 $X=79655 $Y=82290 $D=1
M11 130 129 207 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=79845 $Y=82290 $D=1
M12 208 129 130 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80035 $Y=82290 $D=1
M13 37 131 208 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80225 $Y=82290 $D=1
M14 209 131 37 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80415 $Y=82290 $D=1
M15 130 129 209 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80605 $Y=82290 $D=1
M16 210 129 130 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80795 $Y=82290 $D=1
M17 37 131 210 211 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.27e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=80985 $Y=82290 $D=1
M18 40 130 37 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=4.27e-14 PD=6.7e-07 PS=1.11e-06 $X=81175 $Y=82290 $D=1
M19 37 130 40 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=81365 $Y=82290 $D=1
M20 40 130 37 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=81555 $Y=82290 $D=1
M21 37 130 40 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=81745 $Y=82290 $D=1
M22 40 130 37 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=81935 $Y=82290 $D=1
M23 37 130 40 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=82125 $Y=82290 $D=1
M24 40 130 37 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.73e-14 AS=2.73e-14 PD=6.7e-07 PS=6.7e-07 $X=82315 $Y=82290 $D=1
M25 37 130 40 211 NMOS_VTL L=5e-08 W=1.95e-07 AD=2.0475e-14 AS=2.73e-14 PD=6e-07 PS=6.7e-07 $X=82505 $Y=82290 $D=1
M26 202 37 124 213 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=77360 $Y=83195 $D=0
M27 28 125 202 213 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=77550 $Y=83195 $D=0
M28 28 128 126 213 PMOS_VTL L=5e-08 W=3.15e-07 AD=5.145e-14 AS=3.3075e-14 PD=1.12e-06 PS=8.4e-07 $X=77890 $Y=83195 $D=0
M29 203 124 28 213 PMOS_VTL L=5e-08 W=4.2e-07 AD=5.88e-14 AS=5.145e-14 PD=1.12e-06 PS=1.12e-06 $X=78080 $Y=83090 $D=0
M30 129 126 203 213 PMOS_VTL L=5e-08 W=4.2e-07 AD=4.245e-14 AS=5.88e-14 PD=1.16e-06 PS=1.12e-06 $X=78270 $Y=83090 $D=0
M31 204 128 129 213 PMOS_VTL L=5e-08 W=9e-08 AD=1.26e-14 AS=4.245e-14 PD=4.6e-07 PS=1.16e-06 $X=78480 $Y=83280 $D=0
M32 28 127 204 213 PMOS_VTL L=5e-08 W=9e-08 AD=5.085e-14 AS=1.26e-14 PD=1.55e-06 PS=4.6e-07 $X=78670 $Y=83280 $D=0
M33 127 129 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=5.085e-14 PD=1.54e-06 PS=1.55e-06 $X=78865 $Y=82880 $D=0
M34 28 129 127 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=79055 $Y=82880 $D=0
M35 28 131 128 213 PMOS_VTL L=5e-08 W=3.15e-07 AD=8.19e-14 AS=5.04e-14 PD=1.57e-06 PS=9.5e-07 $X=79450 $Y=82990 $D=0
M36 130 131 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.19e-14 PD=1.54e-06 PS=1.57e-06 $X=79655 $Y=82880 $D=0
M37 28 129 130 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=79845 $Y=82880 $D=0
M38 130 129 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80035 $Y=82880 $D=0
M39 28 131 130 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80225 $Y=82880 $D=0
M40 130 131 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80415 $Y=82880 $D=0
M41 28 129 130 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80605 $Y=82880 $D=0
M42 130 129 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80795 $Y=82880 $D=0
M43 28 131 130 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=80985 $Y=82880 $D=0
M44 40 130 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=81175 $Y=82880 $D=0
M45 28 130 40 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=81365 $Y=82880 $D=0
M46 40 130 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=81555 $Y=82880 $D=0
M47 28 130 40 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=81745 $Y=82880 $D=0
M48 40 130 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=81935 $Y=82880 $D=0
M49 28 130 40 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=82125 $Y=82880 $D=0
M50 40 130 28 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=82315 $Y=82880 $D=0
M51 28 130 40 213 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=82505 $Y=82880 $D=0
X694 27 37 28 24 212 213 CLKBUF_X3 $T=83840 85000 1 0 $X=83725 $Y=83485
X962 164 1 37 28 54 98 214 DFF_X1 $T=1000 79400 0 0 $X=885 $Y=79285
X963 132 1 37 28 41 211 214 DFF_X1 $T=1000 82200 1 0 $X=885 $Y=80685
X964 165 1 37 28 60 212 213 DFF_X1 $T=1000 85000 1 0 $X=885 $Y=83485
X965 166 1 37 28 61 212 213 DFF_X1 $T=4230 85000 1 0 $X=4115 $Y=83485
X966 182 1 37 28 62 211 213 DFF_X1 $T=6700 82200 0 0 $X=6585 $Y=82085
X967 167 1 37 28 29 211 214 DFF_X1 $T=11450 82200 1 0 $X=11335 $Y=80685
X968 168 1 37 28 63 212 213 DFF_X1 $T=11830 85000 1 0 $X=11715 $Y=83485
X969 169 1 37 28 43 212 213 DFF_X1 $T=15060 85000 1 0 $X=14945 $Y=83485
X970 183 1 37 28 30 211 214 DFF_X1 $T=20950 82200 0 180 $X=17605 $Y=80685
X971 106 1 37 28 31 212 213 DFF_X1 $T=18290 85000 1 0 $X=18175 $Y=83485
X972 184 1 37 28 64 211 214 DFF_X1 $T=24180 82200 0 180 $X=20835 $Y=80685
X973 170 1 37 28 32 212 213 DFF_X1 $T=21520 85000 1 0 $X=21405 $Y=83485
X974 136 1 37 28 65 211 213 DFF_X1 $T=27600 82200 0 0 $X=27485 $Y=82085
X975 171 7 37 28 45 211 214 DFF_X1 $T=30450 82200 1 0 $X=30335 $Y=80685
X976 172 1 37 28 46 212 213 DFF_X1 $T=31210 85000 1 0 $X=31095 $Y=83485
X977 173 7 37 28 48 98 214 DFF_X1 $T=34440 79400 0 0 $X=34325 $Y=79285
X978 185 7 37 28 55 212 213 DFF_X1 $T=40140 85000 0 180 $X=36795 $Y=83485
X979 174 7 37 28 56 211 214 DFF_X1 $T=43180 82200 1 0 $X=43065 $Y=80685
X980 175 1 37 28 35 212 213 DFF_X1 $T=43180 85000 1 0 $X=43065 $Y=83485
X981 147 1 37 28 66 212 213 DFF_X1 $T=48120 85000 1 0 $X=48005 $Y=83485
X982 176 1 37 28 67 212 213 DFF_X1 $T=56290 85000 1 0 $X=56175 $Y=83485
X983 177 1 37 28 51 212 213 DFF_X1 $T=59520 85000 1 0 $X=59405 $Y=83485
X984 178 1 37 28 38 211 213 DFF_X1 $T=62750 82200 0 0 $X=62635 $Y=82085
X985 179 1 37 28 68 212 213 DFF_X1 $T=65980 85000 1 0 $X=65865 $Y=83485
X986 163 1 37 28 58 98 214 DFF_X1 $T=74720 79400 0 0 $X=74605 $Y=79285
X987 180 1 37 28 52 212 213 DFF_X1 $T=74720 85000 1 0 $X=74605 $Y=83485
X988 181 1 37 28 59 212 213 DFF_X1 $T=80610 85000 1 0 $X=80495 $Y=83485
X989 162 1 37 28 53 211 214 DFF_X1 $T=81560 82200 1 0 $X=81445 $Y=80685
X1109 194 37 28 69 211 213 CLKBUF_X1 $T=33680 82200 1 180 $X=32995 $Y=82085
X1110 138 37 28 171 212 213 CLKBUF_X1 $T=35770 85000 0 180 $X=35085 $Y=83485
X1111 195 37 28 88 211 213 CLKBUF_X1 $T=36530 82200 1 180 $X=35845 $Y=82085
X1112 140 37 28 173 211 213 CLKBUF_X1 $T=38430 82200 1 180 $X=37745 $Y=82085
X1113 141 37 28 34 211 214 CLKBUF_X1 $T=39000 82200 0 180 $X=38315 $Y=80685
X1114 143 37 28 49 211 214 CLKBUF_X1 $T=41090 82200 0 180 $X=40405 $Y=80685
X1115 142 37 28 185 212 213 CLKBUF_X1 $T=41470 85000 0 180 $X=40785 $Y=83485
X1116 145 37 28 174 212 213 CLKBUF_X1 $T=42610 85000 1 0 $X=42495 $Y=83485
X1117 24 37 28 131 212 213 CLKBUF_X1 $T=79660 85000 1 0 $X=79545 $Y=83485
X1225 39 26 37 28 125 211 214 OR2_X1 $T=73770 82200 1 0 $X=73655 $Y=80685
X1226 39 26 37 28 73 98 214 OR2_X1 $T=73960 79400 0 0 $X=73845 $Y=79285
X1227 39 26 37 28 116 212 213 OR2_X1 $T=77950 85000 1 0 $X=77835 $Y=83485
X1310 36 2 37 28 164 98 214 AND2_X1 $T=5750 79400 0 0 $X=5635 $Y=79285
X1311 36 99 37 28 132 211 214 AND2_X1 $T=6700 82200 0 180 $X=5825 $Y=80685
X1312 36 100 37 28 165 211 213 AND2_X1 $T=6700 82200 1 180 $X=5825 $Y=82085
X1313 36 101 37 28 166 211 214 AND2_X1 $T=6700 82200 1 0 $X=6585 $Y=80685
X1314 36 102 37 28 182 211 214 AND2_X1 $T=11450 82200 0 180 $X=10575 $Y=80685
X1315 36 103 37 28 168 98 214 AND2_X1 $T=12020 79400 0 0 $X=11905 $Y=79285
X1316 36 104 37 28 167 98 214 AND2_X1 $T=15060 79400 0 0 $X=14945 $Y=79285
X1317 36 105 37 28 169 211 214 AND2_X1 $T=17720 82200 0 180 $X=16845 $Y=80685
X1318 36 107 37 28 183 98 214 AND2_X1 $T=20190 79400 1 180 $X=19315 $Y=79285
X1319 36 4 37 28 106 98 214 AND2_X1 $T=20950 79400 0 0 $X=20835 $Y=79285
X1320 36 5 37 28 184 98 214 AND2_X1 $T=23610 79400 1 180 $X=22735 $Y=79285
X1321 36 108 37 28 170 98 214 AND2_X1 $T=26080 79400 0 0 $X=25965 $Y=79285
X1322 36 109 37 28 136 211 214 AND2_X1 $T=28930 82200 0 180 $X=28055 $Y=80685
X1323 36 110 37 28 172 211 214 AND2_X1 $T=29690 82200 1 0 $X=29575 $Y=80685
X1324 47 8 37 28 194 211 213 AND2_X1 $T=34440 82200 1 180 $X=33565 $Y=82085
X1325 47 9 37 28 138 212 213 AND2_X1 $T=35200 85000 0 180 $X=34325 $Y=83485
X1326 47 10 37 28 195 212 213 AND2_X1 $T=35770 85000 1 0 $X=35655 $Y=83485
X1327 47 11 37 28 140 211 213 AND2_X1 $T=37100 82200 0 0 $X=36985 $Y=82085
X1328 47 12 37 28 141 211 214 AND2_X1 $T=39760 82200 0 180 $X=38885 $Y=80685
X1329 47 13 37 28 143 211 214 AND2_X1 $T=39760 82200 1 0 $X=39645 $Y=80685
X1330 36 111 37 28 175 211 213 AND2_X1 $T=40140 82200 0 0 $X=40025 $Y=82085
X1331 47 14 37 28 142 212 213 AND2_X1 $T=40900 85000 0 180 $X=40025 $Y=83485
X1332 47 15 37 28 145 212 213 AND2_X1 $T=41850 85000 1 0 $X=41735 $Y=83485
X1333 36 112 37 28 147 212 213 AND2_X1 $T=46410 85000 1 0 $X=46295 $Y=83485
X1334 36 113 37 28 176 211 213 AND2_X1 $T=52680 82200 1 180 $X=51805 $Y=82085
X1335 36 114 37 28 177 211 213 AND2_X1 $T=52680 82200 0 0 $X=52565 $Y=82085
X1336 36 115 37 28 178 211 213 AND2_X1 $T=61040 82200 0 0 $X=60925 $Y=82085
X1337 36 117 37 28 179 211 213 AND2_X1 $T=65980 82200 0 0 $X=65865 $Y=82085
X1338 36 118 37 28 180 211 213 AND2_X1 $T=66930 82200 0 0 $X=66815 $Y=82085
X1339 36 119 37 28 181 211 213 AND2_X1 $T=71870 82200 0 0 $X=71755 $Y=82085
X1340 36 120 37 28 162 211 214 AND2_X1 $T=73010 82200 0 180 $X=72135 $Y=80685
X1341 36 121 37 28 163 211 214 AND2_X1 $T=73010 82200 1 0 $X=72895 $Y=80685
X1342 36 122 37 28 90 98 214 AND2_X1 $T=73200 79400 0 0 $X=73085 $Y=79285
X1353 186 3 99 42 37 28 98 214 OAI21_X1 $T=8220 79400 0 0 $X=8105 $Y=79285
X1354 133 3 100 42 37 28 211 214 OAI21_X1 $T=8410 82200 1 0 $X=8295 $Y=80685
X1355 134 3 101 42 37 28 211 214 OAI21_X1 $T=9930 82200 0 180 $X=9055 $Y=80685
X1356 198 3 102 42 37 28 98 214 OAI21_X1 $T=11260 79400 0 0 $X=11145 $Y=79285
X1357 78 3 103 42 37 28 98 214 OAI21_X1 $T=13920 79400 1 180 $X=13045 $Y=79285
X1358 79 3 104 42 37 28 98 214 OAI21_X1 $T=16580 79400 0 0 $X=16465 $Y=79285
X1359 80 3 105 42 37 28 98 214 OAI21_X1 $T=18100 79400 1 180 $X=17225 $Y=79285
X1360 81 3 107 42 37 28 98 214 OAI21_X1 $T=20950 79400 1 180 $X=20075 $Y=79285
X1361 82 6 108 44 37 28 98 214 OAI21_X1 $T=25320 79400 0 0 $X=25205 $Y=79285
X1362 135 6 109 44 37 28 211 214 OAI21_X1 $T=27410 82200 1 0 $X=27295 $Y=80685
X1363 137 6 110 44 37 28 98 214 OAI21_X1 $T=29690 79400 1 180 $X=28815 $Y=79285
X1364 139 6 111 44 37 28 211 214 OAI21_X1 $T=36530 82200 1 0 $X=36415 $Y=80685
X1365 144 6 112 44 37 28 211 214 OAI21_X1 $T=41660 82200 1 0 $X=41545 $Y=80685
X1366 146 6 113 44 37 28 211 213 OAI21_X1 $T=47550 82200 0 0 $X=47435 $Y=82085
X1367 196 6 114 44 37 28 211 213 OAI21_X1 $T=50400 82200 1 180 $X=49525 $Y=82085
X1368 197 6 115 44 37 28 211 213 OAI21_X1 $T=55340 82200 0 0 $X=55225 $Y=82085
X1369 200 6 117 44 37 28 211 213 OAI21_X1 $T=58570 82200 0 0 $X=58455 $Y=82085
X1370 152 6 118 44 37 28 211 214 OAI21_X1 $T=63130 82200 1 0 $X=63015 $Y=80685
X1371 156 6 119 44 37 28 211 213 OAI21_X1 $T=67690 82200 0 0 $X=67575 $Y=82085
X1372 123 6 120 44 37 28 211 214 OAI21_X1 $T=69020 82200 0 180 $X=68145 $Y=80685
X1373 201 6 122 44 37 28 98 214 OAI21_X1 $T=69970 79400 0 0 $X=69855 $Y=79285
X1374 160 6 121 44 37 28 211 214 OAI21_X1 $T=69970 82200 1 0 $X=69855 $Y=80685
X1375 158 6 72 44 37 28 98 214 OAI21_X1 $T=71490 79400 0 0 $X=71375 $Y=79285
X1376 74 37 28 186 98 214 INV_X1 $T=7840 79400 0 0 $X=7725 $Y=79285
X1377 75 37 28 133 98 214 INV_X1 $T=9360 79400 1 180 $X=8865 $Y=79285
X1378 76 37 28 134 98 214 INV_X1 $T=10500 79400 1 180 $X=10005 $Y=79285
X1379 77 37 28 198 98 214 INV_X1 $T=13160 79400 1 180 $X=12665 $Y=79285
X1380 83 37 28 135 98 214 INV_X1 $T=26840 79400 0 0 $X=26725 $Y=79285
X1381 84 37 28 137 98 214 INV_X1 $T=28550 79400 0 0 $X=28435 $Y=79285
X1382 85 37 28 139 98 214 INV_X1 $T=32160 79400 0 0 $X=32045 $Y=79285
X1383 86 37 28 144 98 214 INV_X1 $T=37670 79400 0 0 $X=37555 $Y=79285
X1384 26 37 28 47 211 214 INV_X1 $T=41090 82200 1 0 $X=40975 $Y=80685
X1385 87 37 28 146 98 214 INV_X1 $T=42800 79400 0 0 $X=42685 $Y=79285
X1386 50 37 28 196 211 214 INV_X1 $T=46410 82200 1 0 $X=46295 $Y=80685
X1387 148 37 28 197 211 214 INV_X1 $T=49260 82200 1 0 $X=49145 $Y=80685
X1388 150 37 28 200 211 214 INV_X1 $T=51920 82200 1 0 $X=51805 $Y=80685
X1389 149 37 28 152 211 214 INV_X1 $T=56480 82200 1 0 $X=56365 $Y=80685
X1390 153 37 28 123 211 214 INV_X1 $T=58760 82200 1 0 $X=58645 $Y=80685
X1391 190 37 28 156 211 214 INV_X1 $T=61610 82200 1 0 $X=61495 $Y=80685
X1392 157 37 28 158 211 214 INV_X1 $T=61990 82200 1 0 $X=61875 $Y=80685
X1393 154 37 28 201 211 214 INV_X1 $T=64650 82200 1 0 $X=64535 $Y=80685
X1394 159 37 28 160 211 214 INV_X1 $T=66550 82200 1 0 $X=66435 $Y=80685
X1395 161 37 28 57 98 214 INV_X1 $T=69590 79400 0 0 $X=69475 $Y=79285
X1396 26 37 28 36 211 213 INV_X1 $T=70160 82200 0 0 $X=70045 $Y=82085
X1404 148 187 16 37 28 70 98 214 HA_X1 $T=47930 79400 1 180 $X=45915 $Y=79285
X1405 150 188 17 37 28 187 98 214 HA_X1 $T=49830 79400 1 180 $X=47815 $Y=79285
X1406 149 189 18 37 28 188 98 214 HA_X1 $T=51730 79400 1 180 $X=49715 $Y=79285
X1407 153 199 19 37 28 189 98 214 HA_X1 $T=53630 79400 1 180 $X=51615 $Y=79285
X1408 190 151 20 37 28 199 98 214 HA_X1 $T=55530 79400 1 180 $X=53515 $Y=79285
X1409 157 191 21 37 28 151 98 214 HA_X1 $T=57430 79400 1 180 $X=55415 $Y=79285
X1410 154 155 91 37 28 191 211 214 HA_X1 $T=59710 82200 1 0 $X=59595 $Y=80685
X1411 159 192 22 37 28 155 98 214 HA_X1 $T=63320 79400 1 180 $X=61305 $Y=79285
X1412 71 193 23 37 28 192 98 214 HA_X1 $T=65220 79400 1 180 $X=63205 $Y=79285
X1413 161 89 25 37 28 193 98 214 HA_X1 $T=67120 79400 1 180 $X=65105 $Y=79285
X1420 37 116 24 28 37 1 212 213 CLKGATETST_X1 $T=62940 85000 1 0 $X=62825 $Y=83485
.ENDS
***************************************
.SUBCKT ICV_7
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT NOR2_X1 A2 VDD A1 ZN VSS 6 7
** N=8 EP=7 IP=0 FDC=4
M0 ZN A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A1 ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 8 A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 ZN A1 8 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XNOR2_X1 VSS A ZN B VDD 6 7
** N=11 EP=7 IP=0 FDC=10
M0 11 A 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=155 $Y=90 $D=1
M1 VSS B 11 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=345 $Y=90 $D=1
M2 9 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=540 $Y=90 $D=1
M3 ZN A 9 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 9 B ZN 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=920 $Y=90 $D=1
M5 8 A VDD 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=155 $Y=995 $D=0
M6 VDD B 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=345 $Y=995 $D=0
M7 ZN 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=540 $Y=680 $D=0
M8 10 A ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
M9 VDD B 10 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=920 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT XOR2_X1 VDD A Z B VSS 6 7
** N=11 EP=7 IP=0 FDC=10
M0 8 A VSS 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS B 8 6 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.48e-14 AS=2.94e-14 PD=1.12e-06 PS=7e-07 $X=335 $Y=90 $D=1
M2 Z 8 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.48e-14 PD=1.11e-06 PS=1.12e-06 $X=530 $Y=90 $D=1
M3 11 A Z 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=720 $Y=90 $D=1
M4 VSS B 11 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=910 $Y=90 $D=1
M5 10 A 8 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD B 10 7 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.7725e-14 AS=4.41e-14 PD=1.55e-06 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 9 8 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.7725e-14 PD=1.54e-06 PS=1.55e-06 $X=530 $Y=680 $D=0
M8 Z A 9 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=720 $Y=680 $D=0
M9 9 B Z 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=910 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MUX2_X1 A S B VSS VDD Z 7 8
** N=14 EP=8 IP=0 FDC=12
M0 VSS S 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 13 A VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 10 9 13 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 14 S 10 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=715 $Y=90 $D=1
M4 VSS B 14 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=905 $Y=90 $D=1
M5 Z 10 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=1095 $Y=90 $D=1
M6 VDD S 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M7 11 A VDD 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M8 10 S 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M9 12 9 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=715 $Y=995 $D=0
M10 VDD B 12 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=905 $Y=995 $D=0
M11 Z 10 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=1095 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND2_X1 A2 VSS A1 ZN VDD 6 7
** N=8 EP=7 IP=0 FDC=4
M0 8 A2 VSS 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 ZN A1 8 6 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A2 VDD 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A1 ZN 7 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI21_X1 B2 B1 ZN A VSS VDD 7 8
** N=10 EP=8 IP=0 FDC=6
M0 10 B2 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=185 $Y=90 $D=1
M1 ZN B1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=375 $Y=90 $D=1
M2 VSS A ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=565 $Y=90 $D=1
M3 ZN B2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=185 $Y=680 $D=0
M4 9 B1 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=375 $Y=680 $D=0
M5 VDD A 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=565 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_2x1_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NAND3_X1 A3 VSS A2 A1 VDD ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 9 A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 10 A2 9 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 10 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 VDD A2 ZN 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT AOI221_X1 B2 B1 VDD A C2 VSS C1 ZN 9 10
** N=14 EP=10 IP=0 FDC=10
M0 13 B2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 ZN B1 13 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 VSS A ZN 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 14 C2 VSS 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN C1 14 9 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 VDD B2 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M6 11 B1 VDD 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M7 12 A 11 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M8 ZN C2 12 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
M9 12 C1 ZN 10 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT FA_X1 CO CI B A VDD VSS S 8 9
** N=21 EP=9 IP=0 FDC=28
M0 VSS 10 CO 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.375e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=170 $Y=90 $D=1
M1 19 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=4.375e-14 PD=7e-07 PS=1.11e-06 $X=360 $Y=215 $D=1
M2 10 A 19 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=550 $Y=215 $D=1
M3 11 CI 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.045e-14 AS=2.94e-14 PD=7.1e-07 PS=7e-07 $X=740 $Y=215 $D=1
M4 VSS A 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.045e-14 PD=7e-07 PS=7.1e-07 $X=935 $Y=215 $D=1
M5 11 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.205e-14 AS=2.94e-14 PD=6.3e-07 PS=7e-07 $X=1125 $Y=215 $D=1
M6 13 B VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=1465 $Y=90 $D=1
M7 VSS CI 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1655 $Y=90 $D=1
M8 13 A VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=1845 $Y=90 $D=1
M9 15 10 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=3.15e-14 AS=2.94e-14 PD=7.2e-07 PS=7e-07 $X=2035 $Y=90 $D=1
M10 20 CI 15 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=3.15e-14 PD=7e-07 PS=7.2e-07 $X=2235 $Y=90 $D=1
M11 21 B 20 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=2425 $Y=90 $D=1
M12 VSS A 21 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=2615 $Y=90 $D=1
M13 S 15 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=2805 $Y=90 $D=1
M14 VDD 10 CO 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=170 $Y=680 $D=0
M15 16 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=6.615e-14 PD=9.1e-07 PS=1.54e-06 $X=360 $Y=870 $D=0
M16 10 A 16 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=550 $Y=870 $D=0
M17 12 CI 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.53e-14 AS=4.41e-14 PD=1.07e-06 PS=9.1e-07 $X=740 $Y=870 $D=0
M18 VDD A 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.53e-14 PD=9.1e-07 PS=1.07e-06 $X=935 $Y=945 $D=0
M19 12 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=3.3075e-14 AS=4.41e-14 PD=8.4e-07 PS=9.1e-07 $X=1125 $Y=945 $D=0
M20 14 B VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=1465 $Y=995 $D=0
M21 VDD CI 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1655 $Y=995 $D=0
M22 14 A VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=1845 $Y=995 $D=0
M23 15 10 14 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.725e-14 AS=4.41e-14 PD=9.3e-07 PS=9.1e-07 $X=2035 $Y=995 $D=0
M24 17 CI 15 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.725e-14 PD=9.1e-07 PS=9.3e-07 $X=2235 $Y=995 $D=0
M25 18 B 17 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=2425 $Y=995 $D=0
M26 VDD A 18 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=2615 $Y=995 $D=0
M27 S 15 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=2805 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OAI22_X1 B2 B1 VSS ZN A1 A2 VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 VSS B2 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 10 B1 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A1 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=540 $Y=90 $D=1
M3 10 A2 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=730 $Y=90 $D=1
M4 11 B2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M5 ZN B1 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
M6 12 A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=540 $Y=680 $D=0
M7 VDD A2 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=730 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NOR3_X1 A3 VDD A2 A1 VSS ZN 7 8
** N=10 EP=8 IP=0 FDC=6
M0 ZN A3 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A2 ZN 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A1 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 9 A3 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M4 10 A2 9 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M5 ZN A1 10 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_8 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 155 156
** N=281 EP=134 IP=2972 FDC=1464
X955 70 19 39 38 250 279 280 DFF_X1 $T=1000 76600 1 0 $X=885 $Y=75085
X956 248 2 39 38 213 156 281 DFF_X1 $T=1000 79400 1 0 $X=885 $Y=77885
X957 71 19 39 38 56 279 281 DFF_X1 $T=32350 76600 0 0 $X=32235 $Y=76485
X958 247 37 39 38 67 279 281 DFF_X1 $T=75670 76600 0 0 $X=75555 $Y=76485
X959 249 37 39 38 73 279 280 DFF_X1 $T=78330 76600 1 0 $X=78215 $Y=75085
X960 239 37 39 38 68 155 280 DFF_X1 $T=81560 73800 0 0 $X=81445 $Y=73685
X961 238 37 39 38 64 279 280 DFF_X1 $T=81560 76600 1 0 $X=81445 $Y=75085
X962 72 37 39 38 69 156 281 DFF_X1 $T=81560 79400 1 0 $X=81445 $Y=77885
X1088 98 39 38 51 155 280 CLKBUF_X1 $T=15250 73800 1 180 $X=14565 $Y=73685
X1089 265 39 38 40 155 280 CLKBUF_X1 $T=18860 73800 0 0 $X=18745 $Y=73685
X1247 62 178 39 38 90 155 280 OR2_X1 $T=51350 73800 1 180 $X=50475 $Y=73685
X1248 243 186 39 38 178 155 280 OR2_X1 $T=54580 73800 0 0 $X=54465 $Y=73685
X1333 81 1 39 38 248 155 280 AND2_X1 $T=1000 73800 0 0 $X=885 $Y=73685
X1334 104 184 39 38 181 155 280 AND2_X1 $T=53820 73800 0 0 $X=53705 $Y=73685
X1335 43 199 39 38 94 155 280 AND2_X1 $T=72820 73800 0 0 $X=72705 $Y=73685
X1336 43 200 39 38 249 279 280 AND2_X1 $T=74530 76600 0 180 $X=73655 $Y=75085
X1337 43 36 39 38 247 156 281 AND2_X1 $T=73770 79400 1 0 $X=73655 $Y=77885
X1338 43 201 39 38 238 279 281 AND2_X1 $T=74910 76600 1 180 $X=74035 $Y=76485
X1339 43 202 39 38 95 155 280 AND2_X1 $T=75100 73800 1 180 $X=74225 $Y=73685
X1340 43 203 39 38 239 279 281 AND2_X1 $T=74910 76600 0 0 $X=74795 $Y=76485
X1341 43 204 39 38 96 155 280 AND2_X1 $T=75100 73800 0 0 $X=74985 $Y=73685
X1355 206 10 76 40 39 38 156 281 OAI21_X1 $T=22090 79400 1 0 $X=21975 $Y=77885
X1356 217 10 53 40 39 38 156 281 OAI21_X1 $T=23610 79400 0 180 $X=22735 $Y=77885
X1357 57 25 82 209 39 38 155 280 OAI21_X1 $T=37100 73800 0 0 $X=36985 $Y=73685
X1358 221 240 167 222 39 38 279 280 OAI21_X1 $T=39000 76600 1 0 $X=38885 $Y=75085
X1359 26 171 209 84 39 38 155 280 OAI21_X1 $T=40520 73800 0 0 $X=40405 $Y=73685
X1360 61 28 176 226 39 38 279 280 OAI21_X1 $T=43560 76600 1 0 $X=43445 $Y=75085
X1361 189 178 225 91 39 38 155 280 OAI21_X1 $T=52110 73800 1 180 $X=51235 $Y=73685
X1362 228 181 183 229 39 38 156 281 OAI21_X1 $T=53630 79400 1 0 $X=53515 $Y=77885
X1363 65 188 232 185 39 38 279 281 OAI21_X1 $T=58190 76600 1 180 $X=57315 $Y=76485
X1364 32 33 275 187 39 38 155 280 OAI21_X1 $T=61800 73800 1 180 $X=60925 $Y=73685
X1365 260 35 198 66 39 38 155 280 OAI21_X1 $T=68450 73800 0 0 $X=68335 $Y=73685
X1366 236 10 200 40 39 38 279 281 OAI21_X1 $T=69210 76600 0 0 $X=69095 $Y=76485
X1367 246 10 199 40 39 38 155 280 OAI21_X1 $T=70920 73800 0 0 $X=70805 $Y=73685
X1368 42 10 203 40 39 38 156 281 OAI21_X1 $T=71300 79400 1 0 $X=71185 $Y=77885
X1369 245 10 202 40 39 38 279 280 OAI21_X1 $T=71490 76600 1 0 $X=71375 $Y=75085
X1370 276 10 201 40 39 38 279 281 OAI21_X1 $T=71490 76600 0 0 $X=71375 $Y=76485
X1371 211 10 204 40 39 38 279 281 OAI21_X1 $T=73010 76600 1 180 $X=72135 $Y=76485
X1372 215 39 38 115 156 281 INV_X1 $T=14870 79400 0 180 $X=14375 $Y=77885
X1373 50 39 38 125 156 281 INV_X1 $T=17910 79400 0 180 $X=17415 $Y=77885
X1374 216 39 38 116 156 281 INV_X1 $T=18290 79400 0 180 $X=17795 $Y=77885
X1375 51 39 38 272 156 281 INV_X1 $T=19050 79400 1 0 $X=18935 $Y=77885
X1376 205 39 38 126 279 281 INV_X1 $T=21330 76600 0 0 $X=21215 $Y=76485
X1377 254 39 38 206 279 281 INV_X1 $T=23040 76600 1 180 $X=22545 $Y=76485
X1378 266 39 38 217 279 281 INV_X1 $T=23420 76600 1 180 $X=22925 $Y=76485
X1379 219 39 38 78 156 281 INV_X1 $T=24750 79400 1 0 $X=24635 $Y=77885
X1380 101 39 38 81 156 281 INV_X1 $T=33680 79400 1 0 $X=33565 $Y=77885
X1381 57 39 38 221 279 280 INV_X1 $T=37480 76600 1 0 $X=37365 $Y=75085
X1382 224 39 38 170 279 280 INV_X1 $T=41090 76600 1 0 $X=40975 $Y=75085
X1383 226 39 38 171 279 280 INV_X1 $T=42230 76600 1 0 $X=42115 $Y=75085
X1384 227 39 38 267 279 281 INV_X1 $T=51540 76600 0 0 $X=51425 $Y=76485
X1385 268 39 38 229 279 281 INV_X1 $T=54960 76600 1 180 $X=54465 $Y=76485
X1386 232 39 38 228 279 281 INV_X1 $T=56100 76600 0 0 $X=55985 $Y=76485
X1387 230 39 38 188 279 280 INV_X1 $T=56480 76600 1 0 $X=56365 $Y=75085
X1388 231 39 38 185 279 280 INV_X1 $T=56860 76600 1 0 $X=56745 $Y=75085
X1389 106 39 38 189 155 280 INV_X1 $T=59520 73800 0 0 $X=59405 $Y=73685
X1390 107 39 38 195 155 280 INV_X1 $T=63700 73800 0 0 $X=63585 $Y=73685
X1391 108 39 38 260 155 280 INV_X1 $T=65790 73800 0 0 $X=65675 $Y=73685
X1392 235 39 38 236 279 281 INV_X1 $T=68830 76600 0 0 $X=68715 $Y=76485
X1393 237 39 38 276 156 281 INV_X1 $T=69590 79400 1 0 $X=69475 $Y=77885
X1394 261 39 38 245 279 281 INV_X1 $T=69970 76600 0 0 $X=69855 $Y=76485
X1395 259 39 38 246 279 280 INV_X1 $T=70160 76600 1 0 $X=70045 $Y=75085
X1396 109 39 38 211 156 281 INV_X1 $T=70350 79400 1 0 $X=70235 $Y=77885
X1397 110 39 38 66 155 280 INV_X1 $T=70920 73800 1 180 $X=70425 $Y=73685
X1415 278 112 5 39 38 270 155 280 HA_X1 $T=8980 73800 1 180 $X=6965 $Y=73685
X1416 214 47 6 39 38 251 279 280 HA_X1 $T=10500 76600 1 0 $X=10385 $Y=75085
X1417 271 114 128 39 38 263 155 280 HA_X1 $T=14300 73800 1 180 $X=12285 $Y=73685
X1418 252 48 129 39 38 264 279 280 HA_X1 $T=16390 76600 0 180 $X=14375 $Y=75085
X1419 219 255 130 39 38 218 279 281 HA_X1 $T=25320 76600 1 180 $X=23305 $Y=76485
X1420 254 218 131 39 38 253 279 280 HA_X1 $T=25510 76600 0 180 $X=23495 $Y=75085
X1421 54 256 11 39 38 255 279 281 HA_X1 $T=27220 76600 1 180 $X=25205 $Y=76485
X1422 79 207 164 39 38 256 279 281 HA_X1 $T=29120 76600 1 180 $X=27105 $Y=76485
X1423 80 208 165 39 38 207 156 281 HA_X1 $T=31780 79400 1 0 $X=31665 $Y=77885
X1424 118 220 166 39 38 208 156 281 HA_X1 $T=37860 79400 0 180 $X=35845 $Y=77885
X1425 85 223 169 39 38 220 156 281 HA_X1 $T=40900 79400 0 180 $X=38885 $Y=77885
X1426 86 60 173 39 38 223 156 281 HA_X1 $T=42800 79400 0 180 $X=40785 $Y=77885
X1427 259 233 195 39 38 234 279 280 HA_X1 $T=63890 76600 1 0 $X=63775 $Y=75085
X1428 237 234 196 39 38 244 156 281 HA_X1 $T=64460 79400 1 0 $X=64345 $Y=77885
X1429 235 244 210 39 38 277 279 281 HA_X1 $T=66360 76600 0 0 $X=66245 $Y=76485
X1430 261 277 197 39 38 124 156 281 HA_X1 $T=68260 79400 0 180 $X=66245 $Y=77885
X1513 269 38 10 44 39 155 280 NOR2_X1 $T=2900 73800 1 180 $X=2215 $Y=73685
X1514 7 38 99 52 39 155 280 NOR2_X1 $T=16960 73800 1 180 $X=16275 $Y=73685
X1515 272 38 52 163 39 279 281 NOR2_X1 $T=19430 76600 0 0 $X=19315 $Y=76485
X1516 58 38 59 240 39 279 280 NOR2_X1 $T=37860 76600 1 0 $X=37745 $Y=75085
X1517 221 38 58 168 39 279 280 NOR2_X1 $T=39000 76600 0 180 $X=38315 $Y=75085
X1518 26 38 59 273 39 279 280 NOR2_X1 $T=39760 76600 1 0 $X=39645 $Y=75085
X1519 257 38 180 227 39 279 281 NOR2_X1 $T=50210 76600 0 0 $X=50095 $Y=76485
X1520 184 38 104 268 39 155 280 NOR2_X1 $T=53250 73800 0 0 $X=53135 $Y=73685
X1521 181 38 268 274 39 279 281 NOR2_X1 $T=54010 76600 0 0 $X=53895 $Y=76485
X1522 105 38 31 231 39 155 280 NOR2_X1 $T=57240 73800 0 0 $X=57125 $Y=73685
X1523 188 38 231 258 39 279 280 NOR2_X1 $T=57240 76600 1 0 $X=57125 $Y=75085
X1524 32 38 33 186 39 155 280 NOR2_X1 $T=60470 73800 1 180 $X=59785 $Y=73685
X1525 35 38 110 262 39 155 280 NOR2_X1 $T=69970 73800 0 0 $X=69855 $Y=73685
X1526 39 212 269 3 38 155 280 XNOR2_X1 $T=4040 73800 1 180 $X=2785 $Y=73685
X1527 39 241 174 167 38 156 281 XNOR2_X1 $T=37860 79400 1 0 $X=37745 $Y=77885
X1528 39 168 175 172 38 279 281 XNOR2_X1 $T=41280 76600 0 0 $X=41165 $Y=76485
X1529 39 225 182 176 38 279 280 XNOR2_X1 $T=47930 76600 1 0 $X=47815 $Y=75085
X1530 39 242 190 183 38 156 281 XNOR2_X1 $T=52490 79400 1 0 $X=52375 $Y=77885
X1531 39 63 194 198 38 155 280 XNOR2_X1 $T=67310 73800 0 0 $X=67195 $Y=73685
X1532 38 213 45 250 39 156 281 XOR2_X1 $T=4230 79400 1 0 $X=4115 $Y=77885
X1533 38 77 266 253 39 155 280 XOR2_X1 $T=24370 73800 1 180 $X=23115 $Y=73685
X1534 38 170 177 273 39 279 281 XOR2_X1 $T=42420 76600 0 0 $X=42305 $Y=76485
X1535 38 228 191 274 39 156 281 XOR2_X1 $T=56290 79400 1 0 $X=56175 $Y=77885
X1536 38 65 193 258 39 279 281 XOR2_X1 $T=58190 76600 0 0 $X=58075 $Y=76485
X1537 38 189 192 275 39 279 280 XOR2_X1 $T=60090 76600 1 0 $X=59975 $Y=75085
X1538 38 260 34 262 39 155 280 XOR2_X1 $T=66170 73800 0 0 $X=66055 $Y=73685
X1539 14 17 13 39 38 164 279 280 MUX2_X1 $T=28170 76600 0 180 $X=26725 $Y=75085
X1540 12 17 14 39 38 165 155 280 MUX2_X1 $T=27030 73800 0 0 $X=26915 $Y=73685
X1541 15 17 16 39 38 169 155 280 MUX2_X1 $T=30070 73800 0 0 $X=29955 $Y=73685
X1542 16 17 12 39 38 166 279 280 MUX2_X1 $T=31590 76600 0 180 $X=30145 $Y=75085
X1543 18 17 15 39 38 173 279 280 MUX2_X1 $T=31590 76600 1 0 $X=31475 $Y=75085
X1544 20 17 18 39 38 55 155 280 MUX2_X1 $T=35010 73800 1 180 $X=33565 $Y=73685
X1545 21 17 20 39 38 117 155 280 MUX2_X1 $T=36340 73800 1 180 $X=34895 $Y=73685
X1546 23 17 21 39 38 83 279 280 MUX2_X1 $T=36150 76600 1 0 $X=36035 $Y=75085
X1547 174 17 29 39 38 127 279 281 MUX2_X1 $T=46600 76600 1 180 $X=45155 $Y=76485
X1548 29 17 23 39 38 88 279 280 MUX2_X1 $T=46600 76600 1 0 $X=46485 $Y=75085
X1549 175 17 174 39 38 87 156 281 MUX2_X1 $T=48310 79400 0 180 $X=46865 $Y=77885
X1550 177 17 175 39 38 89 156 281 MUX2_X1 $T=48310 79400 1 0 $X=48195 $Y=77885
X1551 182 17 177 39 38 92 156 281 MUX2_X1 $T=51160 79400 1 0 $X=51045 $Y=77885
X1552 190 17 182 39 38 123 156 281 MUX2_X1 $T=58760 79400 0 180 $X=57315 $Y=77885
X1553 191 17 190 39 38 93 156 281 MUX2_X1 $T=58760 79400 1 0 $X=58645 $Y=77885
X1554 192 17 193 39 38 210 279 281 MUX2_X1 $T=61800 76600 0 0 $X=61685 $Y=76485
X1555 193 17 191 39 38 197 156 281 MUX2_X1 $T=63130 79400 0 180 $X=61685 $Y=77885
X1556 34 17 194 39 38 233 279 280 MUX2_X1 $T=62560 76600 1 0 $X=62445 $Y=75085
X1557 194 17 192 39 38 196 156 281 MUX2_X1 $T=63130 79400 1 0 $X=63015 $Y=77885
X1558 272 39 52 10 38 156 281 NAND2_X1 $T=20000 79400 0 180 $X=19315 $Y=77885
X1559 61 39 28 226 38 279 281 NAND2_X1 $T=43560 76600 0 0 $X=43445 $Y=76485
X1560 105 39 31 230 38 155 280 NAND2_X1 $T=57240 73800 1 180 $X=56555 $Y=73685
X1561 32 39 33 187 38 155 280 NAND2_X1 $T=60470 73800 0 0 $X=60355 $Y=73685
X1562 22 24 241 25 39 38 155 280 AOI21_X1 $T=36340 73800 0 0 $X=36225 $Y=73685
X1563 257 180 242 227 39 38 279 281 AOI21_X1 $T=50780 76600 0 0 $X=50665 $Y=76485
X1564 230 187 179 243 39 38 279 280 AOI21_X1 $T=55530 76600 0 180 $X=54655 $Y=75085
X1565 189 187 65 186 39 38 155 280 AOI21_X1 $T=57810 73800 0 0 $X=57695 $Y=73685
X1569 224 39 273 57 38 222 279 280 NAND3_X1 $T=41090 76600 0 180 $X=40215 $Y=75085
X1570 185 39 229 267 38 243 279 280 NAND3_X1 $T=54770 76600 0 180 $X=53895 $Y=75085
X1571 7 49 38 163 8 39 99 265 155 280 AOI221_X1 $T=16960 73800 0 0 $X=16845 $Y=73685
X1572 257 180 38 179 181 39 267 91 279 280 AOI221_X1 $T=50780 76600 1 0 $X=50665 $Y=75085
X1573 212 157 111 4 38 39 46 155 280 FA_X1 $T=4040 73800 0 0 $X=3925 $Y=73685
X1574 157 158 132 270 38 39 74 279 280 FA_X1 $T=4230 76600 1 0 $X=4115 $Y=75085
X1575 158 159 278 251 38 39 75 156 281 FA_X1 $T=5370 79400 1 0 $X=5255 $Y=77885
X1576 159 160 214 263 38 39 113 156 281 FA_X1 $T=8410 79400 1 0 $X=8295 $Y=77885
X1577 160 161 271 264 38 39 215 279 281 FA_X1 $T=13350 76600 0 0 $X=13235 $Y=76485
X1578 161 162 252 100 38 39 216 279 281 FA_X1 $T=16390 76600 0 0 $X=16275 $Y=76485
X1579 162 9 133 97 38 39 205 155 280 FA_X1 $T=20190 73800 0 0 $X=20075 $Y=73685
X1580 28 27 121 102 38 39 257 155 280 FA_X1 $T=43370 73800 0 0 $X=43255 $Y=73685
X1581 180 30 122 103 38 39 184 155 280 FA_X1 $T=46410 73800 0 0 $X=46295 $Y=73685
X1582 170 26 39 172 120 119 38 155 280 OAI22_X1 $T=40520 73800 1 180 $X=39455 $Y=73685
X1583 225 171 39 224 28 61 38 279 280 OAI22_X1 $T=42610 76600 1 0 $X=42495 $Y=75085
X1584 59 38 58 25 39 84 155 280 NOR3_X1 $T=38810 73800 0 0 $X=38695 $Y=73685
.ENDS
***************************************
.SUBCKT MGC_via2_1x2_HV
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_9 1 2 3 4 5 6 7 8 9 10 11 12 13 14
** N=14 EP=14 IP=18 FDC=56
X0 1 2 3 4 5 6 7 13 14 FA_X1 $T=0 0 0 0 $X=-115 $Y=-115
X1 8 9 10 11 5 6 12 13 14 FA_X1 $T=3040 0 0 0 $X=2925 $Y=-115
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_1
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT MGC_via1_1x2_VH_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT NOR4_X1 A4 VDD A3 A2 A1 ZN VSS 8 9
** N=12 EP=9 IP=0 FDC=8
M0 ZN A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 VSS A3 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 ZN A2 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 VSS A1 ZN 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 11 A3 10 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 ZN A1 12 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT NAND4_X1 A4 VSS A3 A2 A1 ZN VDD 8 9
** N=12 EP=9 IP=0 FDC=8
M0 10 A4 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=145 $Y=90 $D=1
M1 11 A3 10 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=335 $Y=90 $D=1
M2 12 A2 11 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=525 $Y=90 $D=1
M3 ZN A1 12 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 ZN A4 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=145 $Y=680 $D=0
M5 VDD A3 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=335 $Y=680 $D=0
M6 ZN A2 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=525 $Y=680 $D=0
M7 VDD A1 ZN 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR4_X1 A1 A2 A3 A4 VSS VDD ZN 8 9
** N=13 EP=9 IP=0 FDC=10
M0 10 A1 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 VSS A2 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 10 A3 VSS 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 10 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 11 A1 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 12 A2 11 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 13 A3 12 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 13 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 10 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_10 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220
+ 221 247 248
** N=450 EP=223 IP=4124 FDC=3058
M0 312 311 14 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=14650 $Y=71090 $D=1
M1 14 313 312 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=14840 $Y=71090 $D=1
M2 312 69 14 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15030 $Y=71090 $D=1
M3 71 70 312 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15220 $Y=71090 $D=1
M4 312 314 71 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=15410 $Y=71090 $D=1
M5 71 315 312 444 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=15600 $Y=71090 $D=1
M6 80 45 324 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=51535 $Y=73295 $D=1
M7 324 281 80 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51725 $Y=73295 $D=1
M8 325 282 324 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=51915 $Y=73295 $D=1
M9 14 81 325 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=52105 $Y=73295 $D=1
M10 325 82 14 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=52295 $Y=73295 $D=1
M11 326 83 14 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=61955 $Y=73295 $D=1
M12 14 84 326 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=62145 $Y=73295 $D=1
M13 326 31 327 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=62510 $Y=73295 $D=1
M14 327 49 326 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=62700 $Y=73295 $D=1
M15 85 50 327 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=62890 $Y=73295 $D=1
M16 327 293 85 247 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=63080 $Y=73295 $D=1
M17 435 311 68 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=14650 $Y=71680 $D=0
M18 436 313 435 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=14840 $Y=71680 $D=0
M19 71 69 436 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15030 $Y=71680 $D=0
M20 437 70 71 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15220 $Y=71680 $D=0
M21 438 314 437 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=15410 $Y=71680 $D=0
M22 68 315 438 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=15600 $Y=71680 $D=0
M23 439 45 80 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=51535 $Y=72490 $D=0
M24 68 281 439 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51725 $Y=72490 $D=0
M25 80 282 68 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=51915 $Y=72490 $D=0
M26 440 81 80 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=52105 $Y=72490 $D=0
M27 68 82 440 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=52295 $Y=72490 $D=0
M28 441 83 68 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=61955 $Y=72490 $D=0
M29 85 84 441 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=1.9845e-13 AS=8.82e-14 PD=1.89e-06 PS=1.54e-06 $X=62145 $Y=72490 $D=0
M30 442 31 85 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=1.9845e-13 PD=1.54e-06 PS=1.89e-06 $X=62510 $Y=72490 $D=0
M31 68 49 442 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=62700 $Y=72490 $D=0
M32 443 50 68 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=62890 $Y=72490 $D=0
M33 85 293 443 447 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=63080 $Y=72490 $D=0
X1394 4 5 14 68 250 248 449 DFF_X1 $T=1000 62600 0 0 $X=885 $Y=62485
X1395 379 6 14 68 254 446 450 DFF_X1 $T=1000 68200 0 0 $X=885 $Y=68085
X1396 380 6 14 68 251 444 450 DFF_X1 $T=1000 71000 1 0 $X=885 $Y=69485
X1397 381 6 14 68 23 444 447 DFF_X1 $T=1000 71000 0 0 $X=885 $Y=70885
X1398 115 5 14 68 18 445 448 DFF_X1 $T=3470 65400 0 0 $X=3355 $Y=65285
X1399 249 6 14 68 22 444 450 DFF_X1 $T=4230 71000 1 0 $X=4115 $Y=69485
X1400 11 5 14 68 19 445 449 DFF_X1 $T=4800 65400 1 0 $X=4685 $Y=63885
X1401 12 5 14 68 329 446 448 DFF_X1 $T=5750 68200 1 0 $X=5635 $Y=66685
X1402 382 6 14 68 21 446 450 DFF_X1 $T=8600 68200 0 0 $X=8485 $Y=68085
X1403 116 5 14 68 90 248 449 DFF_X1 $T=8980 62600 0 0 $X=8865 $Y=62485
X1404 252 5 14 68 26 445 448 DFF_X1 $T=9170 65400 0 0 $X=9055 $Y=65285
X1405 253 6 14 68 24 446 448 DFF_X1 $T=9740 68200 1 0 $X=9625 $Y=66685
X1406 383 6 14 68 255 446 450 DFF_X1 $T=11830 68200 0 0 $X=11715 $Y=68085
X1407 257 6 14 68 256 446 450 DFF_X1 $T=15060 68200 0 0 $X=14945 $Y=68085
X1408 117 5 14 68 258 446 448 DFF_X1 $T=16200 68200 1 0 $X=16085 $Y=66685
X1409 118 5 14 68 259 445 448 DFF_X1 $T=17340 65400 0 0 $X=17225 $Y=65285
X1410 119 5 14 68 109 444 450 DFF_X1 $T=29120 71000 1 0 $X=29005 $Y=69485
X1411 120 5 14 68 126 247 447 DFF_X1 $T=29880 73800 1 0 $X=29765 $Y=72285
X1412 121 5 14 68 95 247 447 DFF_X1 $T=33110 73800 1 0 $X=32995 $Y=72285
X1413 122 60 14 68 112 247 447 DFF_X1 $T=73960 73800 1 0 $X=73845 $Y=72285
X1414 123 60 14 68 113 444 450 DFF_X1 $T=81560 71000 1 0 $X=81445 $Y=69485
X1415 124 60 14 68 114 444 447 DFF_X1 $T=81560 71000 0 0 $X=81445 $Y=70885
X1628 328 14 68 87 445 449 CLKBUF_X1 $T=2330 65400 0 180 $X=1645 $Y=63885
X1629 384 14 68 252 248 449 CLKBUF_X1 $T=7650 62600 0 0 $X=7535 $Y=62485
X1834 256 31 14 68 129 247 447 OR2_X1 $T=21710 73800 1 0 $X=21595 $Y=72285
X1835 74 268 14 68 31 446 450 OR2_X1 $T=26460 68200 1 180 $X=25585 $Y=68085
X1836 291 45 14 68 136 444 447 OR2_X1 $T=54200 71000 0 0 $X=54085 $Y=70885
X1837 48 292 14 68 291 444 450 OR2_X1 $T=62180 71000 1 0 $X=62065 $Y=69485
X1992 67 1 14 68 328 445 449 AND2_X1 $T=1000 65400 1 0 $X=885 $Y=63885
X1993 86 2 14 68 380 445 448 AND2_X1 $T=1000 65400 0 0 $X=885 $Y=65285
X1994 86 3 14 68 381 446 448 AND2_X1 $T=1000 68200 1 0 $X=885 $Y=66685
X1995 86 7 14 68 379 445 449 AND2_X1 $T=3090 65400 0 180 $X=2215 $Y=63885
X1996 86 8 14 68 382 445 448 AND2_X1 $T=2710 65400 0 0 $X=2595 $Y=65285
X1997 86 9 14 68 249 445 449 AND2_X1 $T=4040 65400 0 180 $X=3165 $Y=63885
X1998 86 10 14 68 253 445 449 AND2_X1 $T=4040 65400 1 0 $X=3925 $Y=63885
X1999 67 13 14 68 384 248 449 AND2_X1 $T=8220 62600 0 0 $X=8105 $Y=62485
X2000 86 15 14 68 383 445 448 AND2_X1 $T=9170 65400 1 180 $X=8295 $Y=65285
X2001 86 17 14 68 257 446 448 AND2_X1 $T=8980 68200 1 0 $X=8865 $Y=66685
X2002 30 260 14 68 318 445 449 AND2_X1 $T=20760 65400 1 0 $X=20645 $Y=63885
X2003 86 35 14 68 108 444 450 AND2_X1 $T=26460 71000 1 0 $X=26345 $Y=69485
X2004 86 36 14 68 94 247 447 AND2_X1 $T=27220 73800 1 0 $X=27105 $Y=72285
X2005 86 37 14 68 164 445 448 AND2_X1 $T=27600 65400 0 0 $X=27485 $Y=65285
X2006 77 40 14 68 79 247 447 AND2_X1 $T=39760 73800 1 0 $X=39645 $Y=72285
X2007 368 304 14 68 56 247 447 AND2_X1 $T=73200 73800 1 0 $X=73085 $Y=72285
X2040 260 30 377 336 14 68 248 449 OAI21_X1 $T=21520 62600 1 180 $X=20645 $Y=62485
X2041 341 269 268 386 14 68 445 448 OAI21_X1 $T=25700 65400 0 0 $X=25585 $Y=65285
X2042 96 41 81 97 14 68 247 447 OAI21_X1 $T=42610 73800 1 0 $X=42495 $Y=72285
X2043 153 291 138 281 14 68 444 447 OAI21_X1 $T=60470 71000 1 180 $X=59595 $Y=70885
X2044 359 296 53 360 14 68 247 447 OAI21_X1 $T=65410 73800 1 0 $X=65295 $Y=72285
X2045 410 14 68 385 446 450 INV_X1 $T=19810 68200 0 0 $X=19695 $Y=68085
X2046 316 14 68 334 445 448 INV_X1 $T=22470 65400 1 180 $X=21975 $Y=65285
X2047 31 14 68 293 247 447 INV_X1 $T=63700 73800 0 180 $X=63205 $Y=72285
X2048 355 14 68 296 247 447 INV_X1 $T=64460 73800 1 0 $X=64345 $Y=72285
X2049 358 14 68 360 247 447 INV_X1 $T=66170 73800 1 0 $X=66055 $Y=72285
X2050 365 14 68 363 247 447 INV_X1 $T=68640 73800 0 180 $X=68145 $Y=72285
X2081 127 329 251 14 68 176 247 447 HA_X1 $T=9550 73800 0 180 $X=7535 $Y=72285
X2082 128 259 255 14 68 91 444 447 HA_X1 $T=16960 71000 0 0 $X=16845 $Y=70885
X2083 144 332 258 14 68 72 247 447 HA_X1 $T=17530 73800 1 0 $X=17415 $Y=72285
X2084 378 404 302 14 68 185 444 447 HA_X1 $T=70350 71000 0 0 $X=70235 $Y=70885
X2085 304 429 307 14 68 300 444 447 HA_X1 $T=74340 71000 0 0 $X=74225 $Y=70885
X2086 373 308 62 14 68 368 444 447 HA_X1 $T=76240 71000 0 0 $X=76125 $Y=70885
X2112 14 16 20 68 14 6 444 447 CLKGATETST_X1 $T=8600 71000 0 0 $X=8485 $Y=70885
X2197 250 68 254 174 14 247 447 NOR2_X1 $T=5560 73800 0 180 $X=4875 $Y=72285
X2198 88 68 330 89 14 247 447 NOR2_X1 $T=14490 73800 1 0 $X=14375 $Y=72285
X2199 409 68 331 177 14 247 447 NOR2_X1 $T=16010 73800 1 0 $X=15895 $Y=72285
X2200 28 68 27 376 14 248 449 NOR2_X1 $T=18670 62600 0 0 $X=18555 $Y=62485
X2201 376 68 333 336 14 446 448 NOR2_X1 $T=19430 68200 1 0 $X=19315 $Y=66685
X2202 92 68 29 333 14 446 448 NOR2_X1 $T=20570 68200 0 180 $X=19885 $Y=66685
X2203 385 68 376 418 14 446 450 NOR2_X1 $T=20190 68200 0 0 $X=20075 $Y=68085
X2204 260 68 30 317 14 248 449 NOR2_X1 $T=21520 62600 0 0 $X=21405 $Y=62485
X2205 334 68 333 335 14 445 448 NOR2_X1 $T=22090 65400 1 180 $X=21405 $Y=65285
X2206 410 68 317 340 14 445 448 NOR2_X1 $T=22850 65400 0 0 $X=22735 $Y=65285
X2207 318 68 317 339 14 446 448 NOR2_X1 $T=23040 68200 1 0 $X=22925 $Y=66685
X2208 93 68 270 269 14 445 449 NOR2_X1 $T=26270 65400 1 0 $X=26155 $Y=63885
X2209 387 68 421 165 14 444 447 NOR2_X1 $T=33870 71000 0 0 $X=33755 $Y=70885
X2210 149 68 38 166 14 444 447 NOR2_X1 $T=36340 71000 0 0 $X=36225 $Y=70885
X2211 40 68 77 167 14 247 447 NOR2_X1 $T=38430 73800 1 0 $X=38315 $Y=72285
X2212 296 68 358 357 14 247 447 NOR2_X1 $T=64840 73800 1 0 $X=64725 $Y=72285
X2213 373 68 52 358 14 444 447 NOR2_X1 $T=65790 71000 1 180 $X=65105 $Y=70885
X2214 378 68 300 365 14 444 447 NOR2_X1 $T=70350 71000 1 180 $X=69665 $Y=70885
X2215 304 68 368 106 14 247 447 NOR2_X1 $T=73200 73800 0 180 $X=72515 $Y=72285
X2216 14 254 175 250 68 444 447 XNOR2_X1 $T=7270 71000 1 180 $X=6015 $Y=70885
X2217 14 418 266 261 68 444 450 XNOR2_X1 $T=21330 71000 1 0 $X=21215 $Y=69485
X2218 14 256 332 31 68 444 447 XNOR2_X1 $T=21330 71000 0 0 $X=21215 $Y=70885
X2219 14 339 264 262 68 446 450 XNOR2_X1 $T=23420 68200 0 0 $X=23305 $Y=68085
X2220 14 341 265 267 68 445 448 XNOR2_X1 $T=24560 65400 0 0 $X=24445 $Y=65285
X2221 14 74 263 268 68 446 448 XNOR2_X1 $T=26460 68200 0 180 $X=25205 $Y=66685
X2222 68 130 33 335 14 444 450 XOR2_X1 $T=23610 71000 0 180 $X=22355 $Y=69485
X2223 68 359 49 357 14 444 447 XOR2_X1 $T=61610 71000 0 0 $X=61495 $Y=70885
X2224 265 31 263 14 68 131 444 450 MUX2_X1 $T=24940 71000 0 180 $X=23495 $Y=69485
X2225 266 31 264 14 68 73 247 447 MUX2_X1 $T=24940 73800 0 180 $X=23495 $Y=72285
X2226 264 31 265 14 68 178 444 447 MUX2_X1 $T=23800 71000 0 0 $X=23685 $Y=70885
X2227 33 31 266 14 68 132 247 447 MUX2_X1 $T=24940 73800 1 0 $X=24825 $Y=72285
X2228 28 14 27 410 68 248 449 NAND2_X1 $T=19240 62600 0 0 $X=19125 $Y=62485
X2229 92 14 29 316 68 445 449 NAND2_X1 $T=19430 65400 1 0 $X=19315 $Y=63885
X2230 335 14 410 419 68 446 448 NAND2_X1 $T=22470 68200 1 0 $X=22355 $Y=66685
X2231 93 14 270 386 68 445 448 NAND2_X1 $T=27030 65400 0 0 $X=26915 $Y=65285
X2232 387 14 421 179 68 444 447 NAND2_X1 $T=34440 71000 0 0 $X=34325 $Y=70885
X2233 373 14 52 355 68 444 447 NAND2_X1 $T=64650 71000 0 0 $X=64535 $Y=70885
X2234 316 32 338 377 14 68 445 449 AOI21_X1 $T=22660 65400 1 0 $X=22545 $Y=63885
X2235 93 270 267 269 14 68 445 449 AOI21_X1 $T=27600 65400 0 180 $X=26725 $Y=63885
X2236 149 38 282 76 14 68 247 447 AOI21_X1 $T=36340 73800 1 0 $X=36225 $Y=72285
X2237 153 47 359 48 14 68 444 450 AOI21_X1 $T=61420 71000 1 0 $X=61305 $Y=69485
X2238 355 47 298 292 14 68 444 447 AOI21_X1 $T=65790 71000 0 0 $X=65675 $Y=70885
X2239 378 300 184 365 14 68 247 447 AOI21_X1 $T=69400 73800 0 180 $X=68525 $Y=72285
X2242 360 14 171 363 68 292 247 447 NAND3_X1 $T=66550 73800 1 0 $X=66435 $Y=72285
X2243 378 300 68 298 56 14 363 281 444 447 AOI221_X1 $T=66550 71000 0 0 $X=66435 $Y=70885
X2244 270 25 186 201 68 14 260 248 449 FA_X1 $T=15630 62600 0 0 $X=15515 $Y=62485
X2245 107 34 163 203 68 14 342 248 449 FA_X1 $T=25890 62600 0 0 $X=25775 $Y=62485
X2246 38 202 343 146 68 14 387 446 448 FA_X1 $T=26460 68200 1 0 $X=26345 $Y=66685
X2247 344 204 342 205 68 14 420 445 449 FA_X1 $T=30640 65400 0 180 $X=27485 $Y=63885
X2248 343 187 188 147 68 14 319 445 448 FA_X1 $T=28360 65400 0 0 $X=28245 $Y=65285
X2249 421 319 430 148 68 14 40 444 450 FA_X1 $T=35390 71000 0 180 $X=32235 $Y=69485
X2250 77 388 390 189 68 14 96 444 450 FA_X1 $T=35390 71000 1 0 $X=35275 $Y=69485
X2251 430 345 190 320 68 14 388 446 450 FA_X1 $T=35580 68200 0 0 $X=35465 $Y=68085
X2252 423 191 168 151 68 14 276 248 449 FA_X1 $T=40520 62600 0 0 $X=40405 $Y=62485
X2253 422 207 42 322 68 14 391 445 448 FA_X1 $T=42040 65400 0 0 $X=41925 $Y=65285
X2254 277 283 348 432 68 14 396 444 450 FA_X1 $T=53820 71000 0 180 $X=50665 $Y=69485
X2255 414 285 101 361 68 14 353 445 449 FA_X1 $T=55910 65400 0 180 $X=52755 $Y=63885
X2256 350 289 349 397 68 14 352 444 450 FA_X1 $T=58380 71000 1 0 $X=58265 $Y=69485
X2257 279 294 354 401 68 14 400 446 450 FA_X1 $T=64650 68200 1 180 $X=61495 $Y=68085
X2258 361 55 367 200 68 14 140 248 449 FA_X1 $T=67690 62600 1 180 $X=64535 $Y=62485
X2259 289 402 427 371 68 14 299 446 450 FA_X1 $T=64650 68200 0 0 $X=64535 $Y=68085
X2260 433 295 103 415 68 14 362 445 449 FA_X1 $T=64840 65400 1 0 $X=64725 $Y=63885
X2261 366 301 173 216 68 14 303 445 448 FA_X1 $T=68830 65400 0 0 $X=68715 $Y=65285
X2262 371 306 434 364 68 14 405 446 450 FA_X1 $T=75480 68200 1 180 $X=72325 $Y=68085
X2263 406 305 372 157 68 14 369 445 449 FA_X1 $T=73960 65400 1 0 $X=73845 $Y=63885
X2264 306 61 408 158 68 14 310 445 448 FA_X1 $T=75480 65400 0 0 $X=75365 $Y=65285
X2265 307 309 221 219 68 14 308 444 450 FA_X1 $T=78520 71000 1 0 $X=78405 $Y=69485
X2266 370 310 220 159 68 14 309 446 448 FA_X1 $T=78710 68200 1 0 $X=78595 $Y=66685
X2267 305 63 125 66 68 14 407 248 449 FA_X1 $T=81750 62600 0 0 $X=81635 $Y=62485
X2268 372 64 65 160 68 14 375 445 448 FA_X1 $T=81750 65400 0 0 $X=81635 $Y=65285
X2269 374 407 375 161 68 14 408 446 448 FA_X1 $T=81750 68200 1 0 $X=81635 $Y=66685
X2270 130 334 14 261 29 92 68 445 448 OAI22_X1 $T=21520 65400 1 180 $X=20455 $Y=65285
X2271 385 336 14 262 130 419 68 446 450 OAI22_X1 $T=22470 68200 0 0 $X=22355 $Y=68085
X2272 145 68 162 377 14 337 248 449 NOR3_X1 $T=23800 62600 1 180 $X=22925 $Y=62485
X2277 75 271 344 150 68 14 272 271 39 321 206 273 445 449 ICV_9 $T=34060 65400 1 0 $X=33945 $Y=63885
X2278 320 272 389 141 68 14 346 389 273 423 111 275 445 448 ICV_9 $T=35960 65400 0 0 $X=35845 $Y=65285
X2279 345 78 422 110 68 14 133 411 275 424 420 347 446 450 ICV_9 $T=38620 68200 0 0 $X=38505 $Y=68085
X2280 390 274 346 411 68 14 134 274 391 431 192 98 444 447 ICV_9 $T=39000 71000 0 0 $X=38885 $Y=70885
X2281 321 43 99 412 68 14 392 278 208 194 193 323 445 449 ICV_9 $T=43560 65400 1 0 $X=43445 $Y=63885
X2282 431 276 142 398 68 14 393 413 394 425 195 395 446 450 ICV_9 $T=44700 68200 0 0 $X=44585 $Y=68085
X2283 180 277 347 413 68 14 135 181 279 395 393 287 444 447 ICV_9 $T=45080 71000 0 0 $X=44965 $Y=70885
X2284 322 278 100 392 68 14 394 424 280 209 414 348 446 448 ICV_9 $T=45270 68200 1 0 $X=45155 $Y=66685
X2285 432 433 323 196 68 14 397 283 284 426 286 349 446 450 ICV_9 $T=50780 68200 0 0 $X=50665 $Y=68085
X2286 412 44 169 143 68 14 285 288 46 211 197 351 248 449 ICV_9 $T=52490 62600 0 0 $X=52375 $Y=62485
X2287 182 287 350 396 68 14 137 183 290 352 400 139 247 447 ICV_9 $T=55720 73800 1 0 $X=55605 $Y=72285
X2288 398 210 212 399 68 14 426 399 406 102 154 295 445 449 ICV_9 $T=55910 65400 1 0 $X=55795 $Y=63885
X2289 280 288 198 152 68 14 286 425 199 353 213 401 446 448 ICV_9 $T=56480 68200 1 0 $X=56365 $Y=66685
X2290 354 362 356 351 68 14 402 356 54 104 374 364 446 448 ICV_9 $T=62560 68200 1 0 $X=62445 $Y=66685
X2291 284 51 170 403 68 14 427 294 297 215 214 417 445 448 ICV_9 $T=62750 65400 0 0 $X=62635 $Y=65285
X2292 415 57 172 428 68 14 416 367 217 218 155 428 248 449 ICV_9 $T=67690 62600 0 0 $X=67575 $Y=62485
X2293 297 58 105 416 68 14 301 403 59 369 156 434 445 449 ICV_9 $T=67880 65400 1 0 $X=67765 $Y=63885
X2294 290 299 366 417 68 14 404 302 303 370 405 429 444 450 ICV_9 $T=68260 71000 1 0 $X=68145 $Y=69485
X2298 337 68 338 340 318 341 14 445 449 NOR4_X1 $T=23420 65400 1 0 $X=23305 $Y=63885
X2299 19 14 18 329 250 409 68 247 447 NAND4_X1 $T=10500 73800 0 180 $X=9435 $Y=72285
X2300 22 14 23 251 254 88 68 247 447 NAND4_X1 $T=11640 73800 1 0 $X=11525 $Y=72285
X2301 256 14 255 24 21 330 68 247 447 NAND4_X1 $T=14490 73800 0 180 $X=13425 $Y=72285
X2302 258 14 259 26 90 331 68 247 447 NAND4_X1 $T=17530 73800 0 180 $X=16465 $Y=72285
X2303 250 329 18 19 14 68 315 444 450 OR4_X1 $T=9930 71000 1 0 $X=9815 $Y=69485
X2304 251 23 22 21 14 68 311 444 447 OR4_X1 $T=12590 71000 1 180 $X=11335 $Y=70885
X2305 254 24 255 256 14 68 313 444 447 OR4_X1 $T=13350 71000 0 0 $X=13235 $Y=70885
X2306 90 26 259 258 14 68 314 444 447 OR4_X1 $T=16960 71000 1 180 $X=15705 $Y=70885
.ENDS
***************************************
.SUBCKT MGC_via1_2x1_HV_0
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_11 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 32 33 34 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 268 269
** N=345 EP=194 IP=2953 FDC=1520
X664 72 33 32 11 343 345 CLKBUF_X3 $T=18480 59800 1 0 $X=18365 $Y=58285
X985 311 11 33 32 79 343 345 DFF_X1 $T=4230 59800 1 0 $X=4115 $Y=58285
X986 9 11 33 32 73 269 345 DFF_X1 $T=4800 57000 0 0 $X=4685 $Y=56885
X987 312 13 33 32 34 343 344 DFF_X1 $T=5370 59800 0 0 $X=5255 $Y=59685
X1126 314 33 32 81 343 345 CLKBUF_X1 $T=1760 59800 1 0 $X=1645 $Y=58285
X1127 286 33 32 311 269 345 CLKBUF_X1 $T=2520 57000 0 0 $X=2405 $Y=56885
X1128 313 33 32 124 343 344 CLKBUF_X1 $T=3090 59800 1 180 $X=2405 $Y=59685
X1129 287 33 32 82 268 344 CLKBUF_X1 $T=2710 62600 1 0 $X=2595 $Y=61085
X1130 328 33 32 125 343 344 CLKBUF_X1 $T=3850 59800 0 0 $X=3735 $Y=59685
X1131 315 33 32 126 268 344 CLKBUF_X1 $T=4610 62600 1 0 $X=4495 $Y=61085
X1392 127 2 33 32 80 269 345 AND2_X1 $T=1760 57000 1 180 $X=885 $Y=56885
X1393 54 1 33 32 313 343 344 AND2_X1 $T=1000 59800 0 0 $X=885 $Y=59685
X1394 54 3 33 32 286 269 345 AND2_X1 $T=2520 57000 1 180 $X=1645 $Y=56885
X1395 54 4 33 32 314 343 344 AND2_X1 $T=2520 59800 1 180 $X=1645 $Y=59685
X1396 54 5 33 32 287 268 344 AND2_X1 $T=1950 62600 1 0 $X=1835 $Y=61085
X1397 54 6 33 32 328 343 344 AND2_X1 $T=3090 59800 0 0 $X=2975 $Y=59685
X1398 127 7 33 32 83 269 345 AND2_X1 $T=3280 57000 0 0 $X=3165 $Y=56885
X1399 54 8 33 32 128 269 345 AND2_X1 $T=4040 57000 0 0 $X=3925 $Y=56885
X1400 127 70 33 32 312 343 344 AND2_X1 $T=4610 59800 0 0 $X=4495 $Y=59685
X1401 54 10 33 32 315 268 344 AND2_X1 $T=5940 62600 0 180 $X=5065 $Y=61085
X1402 54 12 33 32 55 268 344 AND2_X1 $T=5940 62600 1 0 $X=5825 $Y=61085
X1403 54 16 33 32 84 268 344 AND2_X1 $T=10310 62600 1 0 $X=10195 $Y=61085
X1415 37 20 289 39 33 32 268 344 OAI21_X1 $T=20950 62600 1 0 $X=20835 $Y=61085
X1416 291 33 32 330 343 345 INV_X1 $T=22280 59800 0 180 $X=21785 $Y=58285
X1514 51 32 56 281 33 343 345 NOR2_X1 $T=13160 59800 1 0 $X=13045 $Y=58285
X1515 35 32 56 317 33 343 345 NOR2_X1 $T=15250 59800 0 180 $X=14565 $Y=58285
X1516 45 32 56 318 33 269 345 NOR2_X1 $T=19810 57000 1 180 $X=19125 $Y=56885
X1517 37 32 20 89 33 268 344 NOR2_X1 $T=20380 62600 1 0 $X=20265 $Y=61085
X1518 57 32 38 74 33 269 345 NOR2_X1 $T=21330 57000 0 0 $X=21215 $Y=56885
X1519 330 32 74 290 33 343 344 NOR2_X1 $T=22090 59800 1 180 $X=21405 $Y=59685
X1520 291 32 40 271 33 269 345 NOR2_X1 $T=23040 57000 0 0 $X=22925 $Y=56885
X1521 23 32 40 292 33 343 345 NOR2_X1 $T=24940 59800 0 180 $X=24255 $Y=58285
X1522 59 32 47 134 33 343 344 NOR2_X1 $T=26460 59800 0 0 $X=26345 $Y=59685
X1523 46 32 64 293 33 343 345 NOR2_X1 $T=27030 59800 1 0 $X=26915 $Y=58285
X1524 46 32 48 58 33 343 344 NOR2_X1 $T=27030 59800 0 0 $X=26915 $Y=59685
X1525 49 32 64 135 33 343 344 NOR2_X1 $T=28170 59800 1 180 $X=27485 $Y=59685
X1526 59 32 48 282 33 343 345 NOR2_X1 $T=29120 59800 1 0 $X=29005 $Y=58285
X1527 45 32 60 273 33 268 344 NOR2_X1 $T=29880 62600 1 0 $X=29765 $Y=61085
X1528 51 32 42 319 33 343 345 NOR2_X1 $T=31400 59800 1 0 $X=31285 $Y=58285
X1529 44 32 25 340 33 343 344 NOR2_X1 $T=33870 59800 1 180 $X=33185 $Y=59685
X1530 35 32 62 284 33 343 345 NOR2_X1 $T=36720 59800 1 0 $X=36605 $Y=58285
X1531 35 32 52 294 33 343 344 NOR2_X1 $T=38050 59800 0 0 $X=37935 $Y=59685
X1532 45 32 62 331 33 343 344 NOR2_X1 $T=39190 59800 1 180 $X=38505 $Y=59685
X1533 51 32 60 276 33 343 345 NOR2_X1 $T=39570 59800 1 0 $X=39455 $Y=58285
X1534 46 32 47 277 33 343 344 NOR2_X1 $T=40900 59800 0 0 $X=40785 $Y=59685
X1535 49 32 48 296 33 343 344 NOR2_X1 $T=42990 59800 0 0 $X=42875 $Y=59685
X1536 59 32 25 297 33 343 345 NOR2_X1 $T=43750 59800 0 180 $X=43065 $Y=58285
X1537 44 32 42 295 33 343 345 NOR2_X1 $T=44320 59800 0 180 $X=43635 $Y=58285
X1538 63 32 64 342 33 343 344 NOR2_X1 $T=44890 59800 1 180 $X=44205 $Y=59685
X1539 63 32 48 320 33 343 345 NOR2_X1 $T=45080 59800 1 0 $X=44965 $Y=58285
X1540 44 32 60 278 33 268 344 NOR2_X1 $T=45650 62600 1 0 $X=45535 $Y=61085
X1541 49 32 47 308 33 343 344 NOR2_X1 $T=46220 59800 0 0 $X=46105 $Y=59685
X1542 50 32 64 298 33 343 345 NOR2_X1 $T=49260 59800 0 180 $X=48575 $Y=58285
X1543 46 32 25 336 33 268 344 NOR2_X1 $T=49830 62600 0 180 $X=49145 $Y=61085
X1544 59 32 42 325 33 268 344 NOR2_X1 $T=50400 62600 0 180 $X=49715 $Y=61085
X1545 35 32 69 143 33 343 344 NOR2_X1 $T=50400 59800 0 0 $X=50285 $Y=59685
X1546 45 32 52 65 33 268 344 NOR2_X1 $T=51160 62600 1 0 $X=51045 $Y=61085
X1547 51 32 62 144 33 343 344 NOR2_X1 $T=52110 59800 0 0 $X=51995 $Y=59685
X1548 59 32 60 326 33 343 344 NOR2_X1 $T=52680 59800 0 0 $X=52565 $Y=59685
X1549 46 32 42 337 33 343 344 NOR2_X1 $T=53250 59800 0 0 $X=53135 $Y=59685
X1550 35 32 121 145 33 269 345 NOR2_X1 $T=53630 57000 0 0 $X=53515 $Y=56885
X1551 49 32 25 332 33 343 344 NOR2_X1 $T=53820 59800 0 0 $X=53705 $Y=59685
X1552 45 32 69 341 33 343 345 NOR2_X1 $T=55530 59800 1 0 $X=55415 $Y=58285
X1553 44 32 62 333 33 268 344 NOR2_X1 $T=57050 62600 1 0 $X=56935 $Y=61085
X1554 51 32 52 322 33 343 345 NOR2_X1 $T=57430 59800 1 0 $X=57315 $Y=58285
X1555 63 32 47 309 33 343 344 NOR2_X1 $T=59520 59800 0 0 $X=59405 $Y=59685
X1556 123 32 64 338 33 269 345 NOR2_X1 $T=62750 57000 1 180 $X=62065 $Y=56885
X1557 50 32 48 310 33 343 344 NOR2_X1 $T=62750 59800 1 180 $X=62065 $Y=59685
X1558 51 32 69 279 33 343 345 NOR2_X1 $T=65600 59800 0 180 $X=64915 $Y=58285
X1559 44 32 52 285 33 269 345 NOR2_X1 $T=66740 57000 1 180 $X=66055 $Y=56885
X1560 59 32 62 302 33 343 345 NOR2_X1 $T=67880 59800 0 180 $X=67195 $Y=58285
X1561 50 32 47 280 33 343 344 NOR2_X1 $T=69970 59800 0 0 $X=69855 $Y=59685
X1562 119 32 64 304 33 343 344 NOR2_X1 $T=72060 59800 1 180 $X=71375 $Y=59685
X1563 123 32 48 303 33 343 344 NOR2_X1 $T=73200 59800 1 180 $X=72515 $Y=59685
X1564 46 32 60 104 33 343 344 NOR2_X1 $T=73770 59800 1 180 $X=73085 $Y=59685
X1565 49 32 42 170 33 268 344 NOR2_X1 $T=75100 62600 0 180 $X=74415 $Y=61085
X1566 51 32 121 327 33 343 344 NOR2_X1 $T=74720 59800 0 0 $X=74605 $Y=59685
X1567 63 32 25 106 33 268 344 NOR2_X1 $T=75670 62600 0 180 $X=74985 $Y=61085
X1568 44 32 69 305 33 268 344 NOR2_X1 $T=76620 62600 1 0 $X=76505 $Y=61085
X1569 59 32 52 334 33 343 344 NOR2_X1 $T=77950 59800 0 0 $X=77835 $Y=59685
X1570 46 32 62 155 33 268 344 NOR2_X1 $T=81370 62600 1 0 $X=81255 $Y=61085
X1571 50 32 42 339 33 343 345 NOR2_X1 $T=81560 59800 1 0 $X=81445 $Y=58285
X1572 50 32 25 156 33 343 344 NOR2_X1 $T=81560 59800 0 0 $X=81445 $Y=59685
X1573 49 32 60 157 33 268 344 NOR2_X1 $T=81940 62600 1 0 $X=81825 $Y=61085
X1574 123 32 47 158 33 343 344 NOR2_X1 $T=83270 59800 0 0 $X=83155 $Y=59685
X1575 119 32 47 307 33 343 345 NOR2_X1 $T=84030 59800 0 180 $X=83345 $Y=58285
X1576 63 32 42 159 33 268 344 NOR2_X1 $T=83650 62600 1 0 $X=83535 $Y=61085
X1577 119 32 48 161 33 268 344 NOR2_X1 $T=84220 62600 1 0 $X=84105 $Y=61085
X1578 33 292 164 272 32 343 344 XNOR2_X1 $T=24560 59800 0 0 $X=24445 $Y=59685
X1579 32 36 88 290 33 343 344 XOR2_X1 $T=24560 59800 1 180 $X=23305 $Y=59685
X1580 32 22 133 289 33 268 344 XOR2_X1 $T=24180 62600 1 0 $X=24065 $Y=61085
X1581 57 33 38 291 32 269 345 NAND2_X1 $T=20760 57000 0 0 $X=20645 $Y=56885
X1582 37 33 20 39 32 343 344 NAND2_X1 $T=20950 59800 0 0 $X=20835 $Y=59685
X1583 39 22 163 89 33 32 268 344 AOI21_X1 $T=23420 62600 1 0 $X=23305 $Y=61085
X1588 14 15 288 182 32 33 316 343 345 FA_X1 $T=7460 59800 1 0 $X=7345 $Y=58285
X1589 130 270 34 79 32 33 129 268 344 FA_X1 $T=14110 62600 0 180 $X=10955 $Y=61085
X1590 288 17 281 73 32 33 191 269 345 FA_X1 $T=13160 57000 0 0 $X=13045 $Y=56885
X1591 270 18 317 109 32 33 86 343 344 FA_X1 $T=14870 59800 0 0 $X=14755 $Y=59685
X1592 162 178 318 114 32 33 329 269 345 FA_X1 $T=16200 57000 0 0 $X=16085 $Y=56885
X1593 85 19 316 329 32 33 132 268 344 FA_X1 $T=17340 62600 1 0 $X=17225 $Y=61085
X1594 131 171 183 184 32 33 87 343 344 FA_X1 $T=17910 59800 0 0 $X=17795 $Y=59685
X1595 75 179 282 293 32 33 274 269 345 FA_X1 $T=24560 57000 0 0 $X=24445 $Y=56885
X1596 41 273 319 340 32 33 61 343 344 FA_X1 $T=30260 59800 0 0 $X=30145 $Y=59685
X1597 136 110 283 185 32 33 90 268 344 FA_X1 $T=32920 62600 1 0 $X=32805 $Y=61085
X1598 43 274 172 335 32 33 137 343 345 FA_X1 $T=33680 59800 1 0 $X=33565 $Y=58285
X1599 335 275 186 284 32 33 91 343 344 FA_X1 $T=35010 59800 0 0 $X=34895 $Y=59685
X1600 283 173 187 116 32 33 138 269 345 FA_X1 $T=35390 57000 0 0 $X=35275 $Y=56885
X1601 275 111 294 331 32 33 139 268 344 FA_X1 $T=35960 62600 1 0 $X=35845 $Y=61085
X1602 76 276 295 297 32 33 141 343 345 FA_X1 $T=40140 59800 1 0 $X=40025 $Y=58285
X1603 93 277 296 342 32 33 140 268 344 FA_X1 $T=45650 62600 0 180 $X=42495 $Y=61085
X1604 92 24 174 180 32 33 95 269 345 FA_X1 $T=45460 57000 0 0 $X=45345 $Y=56885
X1605 166 308 320 298 32 33 94 343 345 FA_X1 $T=48690 59800 0 180 $X=45535 $Y=58285
X1606 165 278 325 336 32 33 142 268 344 FA_X1 $T=46220 62600 1 0 $X=46105 $Y=61085
X1607 77 321 299 117 32 33 146 343 345 FA_X1 $T=52490 59800 1 0 $X=52375 $Y=58285
X1608 321 326 337 332 32 33 147 268 344 FA_X1 $T=54010 62600 1 0 $X=53895 $Y=61085
X1609 96 26 175 323 32 33 148 269 345 FA_X1 $T=56100 57000 0 0 $X=55985 $Y=56885
X1610 299 341 322 333 32 33 66 343 344 FA_X1 $T=56480 59800 0 0 $X=56365 $Y=59685
X1611 323 309 310 338 32 33 300 343 345 FA_X1 $T=58950 59800 1 0 $X=58835 $Y=58285
X1612 167 189 193 300 32 33 98 268 344 FA_X1 $T=58950 62600 1 0 $X=58835 $Y=61085
X1613 67 27 149 188 32 33 97 269 345 FA_X1 $T=62180 57000 1 180 $X=59025 $Y=56885
X1614 99 279 285 302 32 33 301 343 345 FA_X1 $T=61990 59800 1 0 $X=61875 $Y=58285
X1615 168 181 150 176 32 33 68 343 344 FA_X1 $T=62750 59800 0 0 $X=62635 $Y=59685
X1616 169 301 177 118 32 33 100 343 344 FA_X1 $T=65790 59800 0 0 $X=65675 $Y=59685
X1617 28 29 53 306 32 33 101 343 345 FA_X1 $T=67880 59800 1 0 $X=67765 $Y=58285
X1618 151 280 303 304 32 33 103 268 344 FA_X1 $T=68830 62600 1 0 $X=68715 $Y=61085
X1619 102 71 112 120 32 33 105 343 345 FA_X1 $T=70920 59800 1 0 $X=70805 $Y=58285
X1620 154 327 305 334 32 33 152 268 344 FA_X1 $T=81370 62600 0 180 $X=78215 $Y=61085
X1621 107 30 324 113 32 33 192 343 344 FA_X1 $T=78520 59800 0 0 $X=78405 $Y=59685
X1622 306 190 153 122 32 33 324 269 345 FA_X1 $T=78710 57000 0 0 $X=78595 $Y=56885
X1623 78 339 160 307 32 33 108 269 345 FA_X1 $T=81750 57000 0 0 $X=81635 $Y=56885
X1624 36 330 33 272 38 57 32 343 345 OAI22_X1 $T=20950 59800 1 0 $X=20835 $Y=58285
X1629 115 32 21 271 23 22 33 269 345 NOR4_X1 $T=23610 57000 0 0 $X=23495 $Y=56885
.ENDS
***************************************
.SUBCKT INV_X2 A ZN VSS VDD 5 6
** N=6 EP=6 IP=0 FDC=4
M0 ZN A VSS 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=160 $Y=90 $D=1
M1 VSS A ZN 5 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=350 $Y=90 $D=1
M2 ZN A VDD 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=160 $Y=680 $D=0
M3 VDD A ZN 6 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=350 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT OR3_X1 A1 A2 A3 VSS VDD ZN 7 8
** N=11 EP=8 IP=0 FDC=8
M0 VSS A1 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 9 A2 VSS 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 VSS A3 9 7 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=525 $Y=90 $D=1
M3 ZN 9 VSS 7 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=715 $Y=90 $D=1
M4 10 A1 9 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M5 11 A2 10 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M6 VDD A3 11 8 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=525 $Y=995 $D=0
M7 ZN 9 VDD 8 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=715 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_12 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 35 36 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 286 287
** N=360 EP=216 IP=2837 FDC=1582
X897 101 3 36 35 63 287 359 DFF_X1 $T=1760 51400 0 0 $X=1645 $Y=51285
X898 305 3 36 35 105 358 360 DFF_X1 $T=1760 54200 0 0 $X=1645 $Y=54085
X899 306 6 36 35 38 358 359 DFF_X1 $T=4420 54200 1 0 $X=4305 $Y=52685
X900 5 3 36 35 64 287 359 DFF_X1 $T=4990 51400 0 0 $X=4875 $Y=51285
X901 7 3 36 35 321 286 360 DFF_X1 $T=5750 57000 1 0 $X=5635 $Y=55485
X902 102 3 36 35 96 358 359 DFF_X1 $T=20760 54200 1 0 $X=20645 $Y=52685
X1035 332 36 35 305 358 359 CLKBUF_X1 $T=1570 54200 1 0 $X=1455 $Y=52685
X1036 322 36 35 306 358 359 CLKBUF_X1 $T=3850 54200 1 0 $X=3735 $Y=52685
X1037 134 36 35 37 286 360 CLKBUF_X1 $T=4610 57000 1 0 $X=4495 $Y=55485
X1303 155 1 36 35 106 287 359 AND2_X1 $T=1000 51400 0 0 $X=885 $Y=51285
X1304 155 2 36 35 332 358 360 AND2_X1 $T=1000 54200 0 0 $X=885 $Y=54085
X1305 93 4 36 35 322 358 359 AND2_X1 $T=3090 54200 1 0 $X=2975 $Y=52685
X1306 156 12 36 35 184 287 359 AND2_X1 $T=20950 51400 0 0 $X=20835 $Y=51285
X1322 315 27 85 86 36 35 358 359 OAI21_X1 $T=61040 54200 1 0 $X=60925 $Y=52685
X1323 309 36 35 308 286 360 INV_X1 $T=24940 57000 0 180 $X=24445 $Y=55485
X1324 319 36 35 97 287 359 INV_X1 $T=25700 51400 1 180 $X=25205 $Y=51285
X1351 315 174 28 36 35 122 358 360 HA_X1 $T=63320 54200 0 0 $X=63205 $Y=54085
X1434 41 35 66 210 36 286 360 NOR2_X1 $T=11450 57000 1 0 $X=11335 $Y=55485
X1435 40 35 67 301 36 358 359 NOR2_X1 $T=13730 54200 0 180 $X=13045 $Y=52685
X1436 40 35 53 94 36 287 359 NOR2_X1 $T=14490 51400 0 0 $X=14375 $Y=51285
X1437 41 35 67 95 36 287 359 NOR2_X1 $T=15060 51400 0 0 $X=14945 $Y=51285
X1438 44 35 66 288 36 358 359 NOR2_X1 $T=16010 54200 1 0 $X=15895 $Y=52685
X1439 90 35 45 318 36 358 360 NOR2_X1 $T=16390 54200 0 0 $X=16275 $Y=54085
X1440 40 35 66 183 36 286 360 NOR2_X1 $T=18100 57000 1 0 $X=17985 $Y=55485
X1441 46 35 11 289 36 286 360 NOR2_X1 $T=19240 57000 1 0 $X=19125 $Y=55485
X1442 12 35 156 68 36 287 359 NOR2_X1 $T=20380 51400 0 0 $X=20265 $Y=51285
X1443 47 35 137 307 36 287 359 NOR2_X1 $T=22660 51400 0 0 $X=22545 $Y=51285
X1444 90 35 139 187 36 286 360 NOR2_X1 $T=27980 57000 0 180 $X=27295 $Y=55485
X1445 69 35 58 293 36 358 359 NOR2_X1 $T=29310 54200 1 0 $X=29195 $Y=52685
X1446 51 35 56 310 36 358 359 NOR2_X1 $T=30450 54200 1 0 $X=30335 $Y=52685
X1447 55 35 53 343 36 287 359 NOR2_X1 $T=35390 51400 0 0 $X=35275 $Y=51285
X1448 76 35 58 295 36 358 359 NOR2_X1 $T=39570 54200 1 0 $X=39455 $Y=52685
X1449 50 35 56 334 36 358 359 NOR2_X1 $T=42040 54200 1 0 $X=41925 $Y=52685
X1450 51 35 54 330 36 358 360 NOR2_X1 $T=42040 54200 0 0 $X=41925 $Y=54085
X1451 51 35 58 296 36 358 360 NOR2_X1 $T=48690 54200 0 0 $X=48575 $Y=54085
X1452 151 35 53 167 36 287 359 NOR2_X1 $T=49070 51400 0 0 $X=48955 $Y=51285
X1453 50 35 54 320 36 358 360 NOR2_X1 $T=50020 54200 0 0 $X=49905 $Y=54085
X1454 82 35 56 325 36 358 359 NOR2_X1 $T=51730 54200 0 180 $X=51045 $Y=52685
X1455 41 35 23 331 36 358 359 NOR2_X1 $T=54390 54200 1 0 $X=54275 $Y=52685
X1456 40 35 148 312 36 287 359 NOR2_X1 $T=54580 51400 0 0 $X=54465 $Y=51285
X1457 50 35 58 297 36 358 360 NOR2_X1 $T=56670 54200 0 0 $X=56555 $Y=54085
X1458 55 35 24 313 36 287 359 NOR2_X1 $T=58380 51400 0 0 $X=58265 $Y=51285
X1459 153 35 56 345 36 287 359 NOR2_X1 $T=58950 51400 0 0 $X=58835 $Y=51285
X1460 82 35 54 314 36 286 360 NOR2_X1 $T=58950 57000 1 0 $X=58835 $Y=55485
X1461 315 35 27 172 36 358 360 NOR2_X1 $T=61420 54200 0 0 $X=61305 $Y=54085
X1462 82 35 58 316 36 286 360 NOR2_X1 $T=65600 57000 1 0 $X=65485 $Y=55485
X1463 88 35 56 336 36 358 359 NOR2_X1 $T=68260 54200 1 0 $X=68145 $Y=52685
X1464 153 35 54 346 36 358 360 NOR2_X1 $T=68830 54200 1 180 $X=68145 $Y=54085
X1465 151 35 24 317 36 287 359 NOR2_X1 $T=69970 51400 0 0 $X=69855 $Y=51285
X1466 55 35 56 299 36 358 359 NOR2_X1 $T=71680 54200 0 180 $X=70995 $Y=52685
X1467 88 35 54 338 36 358 359 NOR2_X1 $T=74150 54200 0 180 $X=73465 $Y=52685
X1468 82 35 152 347 36 358 360 NOR2_X1 $T=73770 54200 0 0 $X=73655 $Y=54085
X1469 153 35 58 348 36 358 360 NOR2_X1 $T=74340 54200 0 0 $X=74225 $Y=54085
X1470 44 35 148 59 36 287 359 NOR2_X1 $T=74530 51400 0 0 $X=74415 $Y=51285
X1471 88 35 58 339 36 358 359 NOR2_X1 $T=75100 54200 1 0 $X=74985 $Y=52685
X1472 153 35 152 349 36 358 359 NOR2_X1 $T=75670 54200 1 0 $X=75555 $Y=52685
X1473 90 35 23 104 36 358 359 NOR2_X1 $T=76240 54200 1 0 $X=76125 $Y=52685
X1474 178 35 112 100 36 287 359 NOR2_X1 $T=77380 51400 0 0 $X=77265 $Y=51285
X1475 82 35 60 300 36 358 359 NOR2_X1 $T=77950 54200 1 0 $X=77835 $Y=52685
X1476 61 35 179 350 36 287 359 NOR2_X1 $T=80800 51400 0 0 $X=80685 $Y=51285
X1477 51 35 91 193 36 286 360 NOR2_X1 $T=82320 57000 1 0 $X=82205 $Y=55485
X1478 180 35 181 356 36 287 359 NOR2_X1 $T=82890 51400 0 0 $X=82775 $Y=51285
X1479 69 35 62 340 36 287 359 NOR2_X1 $T=83460 51400 0 0 $X=83345 $Y=51285
X1480 35 291 186 211 36 358 359 XOR2_X1 $T=25130 54200 0 180 $X=23875 $Y=52685
X1481 35 309 103 351 36 286 360 XOR2_X1 $T=24940 57000 1 0 $X=24825 $Y=55485
X1482 35 319 160 194 36 358 359 XOR2_X1 $T=28170 54200 0 180 $X=26915 $Y=52685
X1483 35 292 49 109 36 287 359 XOR2_X1 $T=31400 51400 0 0 $X=31285 $Y=51285
X1484 46 36 11 290 35 358 360 NAND2_X1 $T=19810 54200 0 0 $X=19695 $Y=54085
X1485 315 36 27 86 35 358 359 NAND2_X1 $T=62370 54200 0 180 $X=61685 $Y=52685
X1486 46 11 351 289 36 35 286 360 AOI21_X1 $T=20570 57000 0 180 $X=19695 $Y=55485
X1487 308 290 185 289 36 35 286 360 AOI21_X1 $T=23800 57000 0 180 $X=22925 $Y=55485
X1488 290 14 212 342 36 35 358 360 AOI21_X1 $T=23230 54200 0 0 $X=23115 $Y=54085
X1489 14 291 309 307 36 35 358 360 AOI21_X1 $T=23990 54200 0 0 $X=23875 $Y=54085
X1490 140 292 319 161 36 35 287 359 AOI21_X1 $T=28360 51400 1 180 $X=27485 $Y=51285
X1495 42 213 321 301 35 36 323 358 360 FA_X1 $T=13350 54200 0 0 $X=13235 $Y=54085
X1496 201 8 323 341 35 36 108 286 360 FA_X1 $T=15060 57000 1 0 $X=14945 $Y=55485
X1497 182 9 324 136 35 36 10 287 359 FA_X1 $T=15630 51400 0 0 $X=15515 $Y=51285
X1498 341 288 318 202 35 36 324 358 359 FA_X1 $T=17720 54200 1 0 $X=17605 $Y=52685
X1499 98 293 162 310 35 36 70 287 359 FA_X1 $T=28360 51400 0 0 $X=28245 $Y=51285
X1500 48 16 203 141 35 36 357 286 360 FA_X1 $T=29120 57000 1 0 $X=29005 $Y=55485
X1501 110 195 214 142 35 36 71 286 360 FA_X1 $T=32160 57000 1 0 $X=32045 $Y=55485
X1502 163 17 164 333 35 36 111 358 360 FA_X1 $T=32350 54200 0 0 $X=32235 $Y=54085
X1503 333 357 196 99 35 36 165 358 360 FA_X1 $T=35390 54200 0 0 $X=35275 $Y=54085
X1504 18 19 343 143 35 36 344 287 359 FA_X1 $T=35960 51400 0 0 $X=35845 $Y=51285
X1505 74 352 77 200 35 36 294 286 360 FA_X1 $T=38620 57000 1 0 $X=38505 $Y=55485
X1506 189 197 344 204 35 36 75 287 359 FA_X1 $T=42040 51400 1 180 $X=38885 $Y=51285
X1507 188 294 79 304 35 36 113 286 360 FA_X1 $T=41660 57000 1 0 $X=41545 $Y=55485
X1508 78 20 205 144 35 36 303 287 359 FA_X1 $T=42040 51400 0 0 $X=41925 $Y=51285
X1509 352 295 330 334 35 36 311 358 360 FA_X1 $T=42610 54200 0 0 $X=42495 $Y=54085
X1510 52 206 80 335 35 36 115 358 359 FA_X1 $T=45080 54200 1 0 $X=44965 $Y=52685
X1511 166 303 207 311 35 36 114 358 360 FA_X1 $T=48690 54200 1 180 $X=45535 $Y=54085
X1512 335 296 320 325 35 36 22 358 359 FA_X1 $T=48120 54200 1 0 $X=48005 $Y=52685
X1513 304 21 81 145 35 36 116 286 360 FA_X1 $T=48690 57000 1 0 $X=48575 $Y=55485
X1514 117 326 83 147 35 36 118 286 360 FA_X1 $T=51730 57000 1 0 $X=51615 $Y=55485
X1515 326 133 312 331 35 36 170 358 359 FA_X1 $T=58000 54200 0 180 $X=54845 $Y=52685
X1516 119 25 313 149 35 36 84 358 359 FA_X1 $T=61040 54200 0 180 $X=57885 $Y=52685
X1517 190 297 314 345 35 36 57 358 360 FA_X1 $T=58380 54200 0 0 $X=58265 $Y=54085
X1518 171 26 173 327 35 36 121 287 359 FA_X1 $T=60850 51400 0 0 $X=60735 $Y=51285
X1519 120 328 87 150 35 36 123 286 360 FA_X1 $T=62560 57000 1 0 $X=62445 $Y=55485
X1520 191 29 198 209 35 36 125 287 359 FA_X1 $T=63890 51400 0 0 $X=63775 $Y=51285
X1521 327 316 346 336 35 36 126 358 360 FA_X1 $T=65220 54200 0 0 $X=65105 $Y=54085
X1522 124 353 298 337 35 36 127 286 360 FA_X1 $T=66170 57000 1 0 $X=66055 $Y=55485
X1523 353 30 175 199 35 36 128 287 359 FA_X1 $T=66930 51400 0 0 $X=66815 $Y=51285
X1524 298 299 176 317 35 36 129 358 360 FA_X1 $T=68830 54200 0 0 $X=68715 $Y=54085
X1525 215 31 177 208 35 36 89 287 359 FA_X1 $T=70540 51400 0 0 $X=70425 $Y=51285
X1526 337 347 348 338 35 36 130 286 360 FA_X1 $T=72440 57000 1 0 $X=72325 $Y=55485
X1527 354 300 349 339 35 36 329 358 360 FA_X1 $T=78710 54200 0 0 $X=78595 $Y=54085
X1528 328 354 32 355 35 36 131 286 360 FA_X1 $T=79280 57000 1 0 $X=79165 $Y=55485
X1529 355 350 356 340 35 36 132 358 359 FA_X1 $T=81750 54200 1 0 $X=81635 $Y=52685
X1530 192 33 329 154 35 36 92 358 360 FA_X1 $T=81750 54200 0 0 $X=81635 $Y=54085
X1531 291 35 307 342 36 158 358 360 NOR3_X1 $T=24750 54200 0 0 $X=24635 $Y=54085
X1532 292 35 161 159 36 302 287 359 NOR3_X1 $T=27600 51400 1 180 $X=26725 $Y=51285
X1533 146 35 168 169 36 292 287 359 NOR3_X1 $T=52110 51400 0 0 $X=51995 $Y=51285
X1542 96 35 64 321 43 107 36 287 359 NOR4_X1 $T=11830 51400 0 0 $X=11715 $Y=51285
X1543 302 35 157 15 138 291 36 287 359 NOR4_X1 $T=24940 51400 1 180 $X=23875 $Y=51285
X1545 135 40 36 35 286 360 INV_X2 $T=8980 57000 1 0 $X=8865 $Y=55485
X1546 39 41 36 35 287 359 INV_X2 $T=9360 51400 0 0 $X=9245 $Y=51285
X1547 321 53 36 35 287 359 INV_X2 $T=10500 51400 1 180 $X=9815 $Y=51285
X1548 65 90 36 35 358 359 INV_X2 $T=11260 54200 1 0 $X=11145 $Y=52685
X1549 63 66 36 35 358 359 INV_X2 $T=11830 54200 1 0 $X=11715 $Y=52685
X1550 43 45 36 35 358 359 INV_X2 $T=13730 54200 1 0 $X=13615 $Y=52685
X1551 38 44 36 35 286 360 INV_X2 $T=18670 57000 1 0 $X=18555 $Y=55485
X1552 141 181 36 35 358 360 INV_X2 $T=30450 54200 0 0 $X=30335 $Y=54085
X1553 72 179 36 35 286 360 INV_X2 $T=35200 57000 1 0 $X=35085 $Y=55485
X1554 73 112 36 35 358 359 INV_X2 $T=37480 54200 1 0 $X=37365 $Y=52685
X1555 68 13 289 36 35 342 286 360 OR3_X1 $T=22090 57000 1 0 $X=21975 $Y=55485
.ENDS
***************************************
.SUBCKT AND4_X1 A1 A2 A3 A4 VSS VDD ZN 8 9
** N=13 EP=9 IP=0 FDC=10
M0 11 A1 10 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.205e-14 PD=7e-07 PS=6.3e-07 $X=145 $Y=90 $D=1
M1 12 A2 11 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=335 $Y=90 $D=1
M2 13 A3 12 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=2.94e-14 AS=2.94e-14 PD=7e-07 PS=7e-07 $X=525 $Y=90 $D=1
M3 VSS A4 13 8 NMOS_VTL L=5e-08 W=2.1e-07 AD=4.375e-14 AS=2.94e-14 PD=1.11e-06 PS=7e-07 $X=715 $Y=90 $D=1
M4 ZN 10 VSS 8 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=4.375e-14 PD=1.04e-06 PS=1.11e-06 $X=905 $Y=90 $D=1
M5 10 A1 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=3.3075e-14 PD=9.1e-07 PS=8.4e-07 $X=145 $Y=995 $D=0
M6 VDD A2 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=335 $Y=995 $D=0
M7 10 A3 VDD 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=4.41e-14 AS=4.41e-14 PD=9.1e-07 PS=9.1e-07 $X=525 $Y=995 $D=0
M8 VDD A4 10 9 PMOS_VTL L=5e-08 W=3.15e-07 AD=6.615e-14 AS=4.41e-14 PD=1.54e-06 PS=9.1e-07 $X=715 $Y=995 $D=0
M9 ZN 10 VDD 9 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=6.615e-14 PD=1.47e-06 PS=1.54e-06 $X=905 $Y=680 $D=0
.ENDS
***************************************
.SUBCKT ICV_13 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 35 36 37 38 39 40 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 58 59 60 61 62 63
+ 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 285 286
** N=362 EP=220 IP=2965 FDC=1578
X1006 311 3 36 35 289 360 361 DFF_X1 $T=1000 48600 0 0 $X=885 $Y=48485
X1007 287 5 36 35 38 286 362 DFF_X1 $T=1760 45800 0 0 $X=1645 $Y=45685
X1008 336 5 36 35 62 285 361 DFF_X1 $T=3850 51400 1 0 $X=3735 $Y=49885
X1009 312 5 36 35 9 360 362 DFF_X1 $T=5560 48600 1 0 $X=5445 $Y=47085
X1010 337 5 36 35 64 286 362 DFF_X1 $T=9170 45800 0 0 $X=9055 $Y=45685
X1011 313 3 36 35 66 360 361 DFF_X1 $T=16960 48600 0 0 $X=16845 $Y=48485
X1012 10 3 36 35 106 286 362 DFF_X1 $T=19050 45800 0 0 $X=18935 $Y=45685
X1135 330 36 35 287 360 362 CLKBUF_X1 $T=1000 48600 1 0 $X=885 $Y=47085
X1136 346 36 35 59 360 362 CLKBUF_X1 $T=1570 48600 1 0 $X=1455 $Y=47085
X1137 134 36 35 60 285 361 CLKBUF_X1 $T=1760 51400 1 0 $X=1645 $Y=49885
X1138 310 36 35 311 285 361 CLKBUF_X1 $T=2900 51400 0 180 $X=2215 $Y=49885
X1139 303 36 35 337 360 362 CLKBUF_X1 $T=3660 48600 1 0 $X=3545 $Y=47085
X1140 288 36 35 312 360 362 CLKBUF_X1 $T=4230 48600 1 0 $X=4115 $Y=47085
X1141 331 36 35 336 360 361 CLKBUF_X1 $T=4230 48600 0 0 $X=4115 $Y=48485
X1142 347 36 35 313 360 362 CLKBUF_X1 $T=11830 48600 1 0 $X=11715 $Y=47085
X1430 58 1 36 35 346 286 362 AND2_X1 $T=1000 45800 0 0 $X=885 $Y=45685
X1431 58 102 36 35 310 285 361 AND2_X1 $T=1000 51400 1 0 $X=885 $Y=49885
X1432 61 2 36 35 330 360 362 AND2_X1 $T=2900 48600 0 180 $X=2025 $Y=47085
X1433 61 4 36 35 303 360 362 AND2_X1 $T=2900 48600 1 0 $X=2785 $Y=47085
X1434 61 6 36 35 331 285 361 AND2_X1 $T=3090 51400 1 0 $X=2975 $Y=49885
X1435 61 7 36 35 288 360 362 AND2_X1 $T=4800 48600 1 0 $X=4685 $Y=47085
X1436 58 8 36 35 347 360 362 AND2_X1 $T=11070 48600 1 0 $X=10955 $Y=47085
X1452 68 13 72 71 36 35 285 361 OAI21_X1 $T=23800 51400 0 180 $X=22925 $Y=49885
X1453 42 19 166 16 36 35 360 361 OAI21_X1 $T=27790 48600 1 180 $X=26915 $Y=48485
X1454 85 25 340 83 36 35 360 362 OAI21_X1 $T=55150 48600 0 180 $X=54275 $Y=47085
X1455 340 36 35 202 360 361 INV_X1 $T=56100 48600 0 0 $X=55985 $Y=48485
X1555 67 35 12 194 36 360 362 NOR2_X1 $T=22090 48600 1 0 $X=21975 $Y=47085
X1556 70 35 12 357 36 360 362 NOR2_X1 $T=23230 48600 0 180 $X=22545 $Y=47085
X1557 69 35 14 305 36 286 362 NOR2_X1 $T=23230 45800 0 0 $X=23115 $Y=45685
X1558 42 35 19 73 36 285 361 NOR2_X1 $T=26840 51400 1 0 $X=26725 $Y=49885
X1559 44 35 142 197 36 285 361 NOR2_X1 $T=29690 51400 1 0 $X=29575 $Y=49885
X1560 76 35 48 198 36 285 361 NOR2_X1 $T=33870 51400 1 0 $X=33755 $Y=49885
X1561 157 35 28 291 36 286 362 NOR2_X1 $T=34820 45800 0 0 $X=34705 $Y=45685
X1562 55 35 77 199 36 285 361 NOR2_X1 $T=36340 51400 1 0 $X=36225 $Y=49885
X1563 45 35 29 317 36 286 362 NOR2_X1 $T=36720 45800 0 0 $X=36605 $Y=45685
X1564 21 35 53 333 36 360 361 NOR2_X1 $T=36910 48600 0 0 $X=36795 $Y=48485
X1565 49 35 78 292 36 360 362 NOR2_X1 $T=39950 48600 1 0 $X=39835 $Y=47085
X1566 79 35 48 47 36 285 361 NOR2_X1 $T=41660 51400 1 0 $X=41545 $Y=49885
X1567 31 35 39 318 36 360 362 NOR2_X1 $T=42040 48600 1 0 $X=41925 $Y=47085
X1568 55 35 145 172 36 285 361 NOR2_X1 $T=44890 51400 0 180 $X=44205 $Y=49885
X1569 49 35 77 200 36 285 361 NOR2_X1 $T=45460 51400 0 180 $X=44775 $Y=49885
X1570 45 35 28 334 36 360 361 NOR2_X1 $T=45080 48600 0 0 $X=44965 $Y=48485
X1571 76 35 53 335 36 360 361 NOR2_X1 $T=46790 48600 0 0 $X=46675 $Y=48485
X1572 55 35 48 294 36 285 361 NOR2_X1 $T=47170 51400 1 0 $X=47055 $Y=49885
X1573 21 35 29 319 36 360 362 NOR2_X1 $T=48120 48600 0 180 $X=47435 $Y=47085
X1574 31 35 77 353 36 360 361 NOR2_X1 $T=49070 48600 0 0 $X=48955 $Y=48485
X1575 21 35 28 295 36 360 361 NOR2_X1 $T=49640 48600 0 0 $X=49525 $Y=48485
X1576 79 35 53 308 36 360 361 NOR2_X1 $T=52490 48600 1 180 $X=51805 $Y=48485
X1577 76 35 29 320 36 360 362 NOR2_X1 $T=53060 48600 0 180 $X=52375 $Y=47085
X1578 83 35 147 54 36 360 362 NOR2_X1 $T=54390 48600 0 180 $X=53705 $Y=47085
X1579 91 35 78 296 36 286 362 NOR2_X1 $T=54010 45800 0 0 $X=53895 $Y=45685
X1580 49 35 48 297 36 360 362 NOR2_X1 $T=56290 48600 1 0 $X=56175 $Y=47085
X1581 76 35 28 118 36 285 361 NOR2_X1 $T=57810 51400 1 0 $X=57695 $Y=49885
X1582 55 35 53 88 36 285 361 NOR2_X1 $T=58380 51400 1 0 $X=58265 $Y=49885
X1583 31 35 145 323 36 360 361 NOR2_X1 $T=58760 48600 0 0 $X=58645 $Y=48485
X1584 93 35 77 329 36 360 361 NOR2_X1 $T=59900 48600 1 180 $X=59215 $Y=48485
X1585 31 35 48 298 36 360 361 NOR2_X1 $T=60850 48600 0 0 $X=60735 $Y=48485
X1586 93 35 145 324 36 360 361 NOR2_X1 $T=61420 48600 0 0 $X=61305 $Y=48485
X1587 91 35 77 325 36 360 362 NOR2_X1 $T=64460 48600 0 180 $X=63775 $Y=47085
X1588 79 35 28 299 36 360 361 NOR2_X1 $T=65220 48600 0 0 $X=65105 $Y=48485
X1589 55 35 29 326 36 360 361 NOR2_X1 $T=65790 48600 0 0 $X=65675 $Y=48485
X1590 49 35 53 354 36 360 361 NOR2_X1 $T=66360 48600 0 0 $X=66245 $Y=48485
X1591 31 35 53 179 36 360 361 NOR2_X1 $T=68070 48600 1 180 $X=67385 $Y=48485
X1592 91 35 145 180 36 360 361 NOR2_X1 $T=68070 48600 0 0 $X=67955 $Y=48485
X1593 93 35 48 204 36 285 361 NOR2_X1 $T=68260 51400 1 0 $X=68145 $Y=49885
X1594 79 35 142 358 36 286 362 NOR2_X1 $T=69400 45800 0 0 $X=69285 $Y=45685
X1595 55 35 182 309 36 286 362 NOR2_X1 $T=71680 45800 1 180 $X=70995 $Y=45685
X1596 49 35 28 342 36 360 362 NOR2_X1 $T=71300 48600 1 0 $X=71185 $Y=47085
X1597 55 35 28 184 36 285 361 NOR2_X1 $T=72060 51400 0 180 $X=71375 $Y=49885
X1598 95 35 150 350 36 360 362 NOR2_X1 $T=73770 48600 0 180 $X=73085 $Y=47085
X1599 44 35 154 302 36 286 362 NOR2_X1 $T=81370 45800 0 0 $X=81255 $Y=45685
X1600 156 35 100 328 36 285 361 NOR2_X1 $T=83270 51400 1 0 $X=83155 $Y=49885
X1601 157 35 56 355 36 286 362 NOR2_X1 $T=83460 45800 0 0 $X=83345 $Y=45685
X1602 36 357 195 290 35 360 361 XNOR2_X1 $T=23800 48600 1 180 $X=22545 $Y=48485
X1603 35 351 103 305 36 360 362 XOR2_X1 $T=26080 48600 0 180 $X=24825 $Y=47085
X1604 35 202 90 121 36 285 361 XOR2_X1 $T=59900 51400 1 0 $X=59785 $Y=49885
X1605 68 36 13 71 35 285 361 NAND2_X1 $T=22470 51400 1 0 $X=22355 $Y=49885
X1606 42 36 19 16 35 360 361 NAND2_X1 $T=24940 48600 0 0 $X=24825 $Y=48485
X1607 17 16 196 104 36 35 285 361 AOI21_X1 $T=24750 51400 1 0 $X=24635 $Y=49885
X1608 140 17 351 15 36 35 360 362 AOI21_X1 $T=26840 48600 0 180 $X=25965 $Y=47085
X1614 314 36 315 65 35 110 360 361 NAND3_X1 $T=16200 48600 0 0 $X=16085 $Y=48485
X1615 141 36 74 316 35 75 286 362 NAND3_X1 $T=28740 45800 0 0 $X=28625 $Y=45685
X1616 191 289 205 138 35 36 111 285 361 FA_X1 $T=14870 51400 1 0 $X=14755 $Y=49885
X1617 193 206 213 137 35 36 40 286 362 FA_X1 $T=19050 45800 1 180 $X=15895 $Y=45685
X1618 192 207 129 128 35 36 112 285 361 FA_X1 $T=17910 51400 1 0 $X=17795 $Y=49885
X1619 18 20 43 332 35 36 113 360 362 FA_X1 $T=26840 48600 1 0 $X=26725 $Y=47085
X1620 332 217 306 216 35 36 170 360 361 FA_X1 $T=33870 48600 0 0 $X=33755 $Y=48485
X1621 306 291 317 333 35 36 114 360 362 FA_X1 $T=36910 48600 1 0 $X=36795 $Y=47085
X1622 46 22 307 352 35 36 115 285 361 FA_X1 $T=38620 51400 1 0 $X=38505 $Y=49885
X1623 352 292 318 130 35 36 171 286 362 FA_X1 $T=40900 45800 0 0 $X=40785 $Y=45685
X1624 307 293 218 348 35 36 173 360 361 FA_X1 $T=42040 48600 0 0 $X=41925 $Y=48485
X1625 293 23 174 131 35 36 116 286 362 FA_X1 $T=44510 45800 0 0 $X=44395 $Y=45685
X1626 348 334 319 335 35 36 50 360 362 FA_X1 $T=44510 48600 1 0 $X=44395 $Y=47085
X1627 51 294 80 353 35 36 321 285 361 FA_X1 $T=48690 51400 1 0 $X=48575 $Y=49885
X1628 52 295 320 308 35 36 339 360 362 FA_X1 $T=49450 48600 1 0 $X=49335 $Y=47085
X1629 201 24 175 146 35 36 338 286 362 FA_X1 $T=54010 45800 1 180 $X=50855 $Y=45685
X1630 84 338 321 339 35 36 81 285 361 FA_X1 $T=54770 51400 0 180 $X=51615 $Y=49885
X1631 322 296 208 148 35 36 176 286 362 FA_X1 $T=57620 45800 1 180 $X=54465 $Y=45685
X1632 117 209 322 349 35 36 87 285 361 FA_X1 $T=54770 51400 1 0 $X=54655 $Y=49885
X1633 86 26 177 149 35 36 119 286 362 FA_X1 $T=57620 45800 0 0 $X=57505 $Y=45685
X1634 349 297 323 329 35 36 120 360 362 FA_X1 $T=57810 48600 1 0 $X=57695 $Y=47085
X1635 89 27 210 221 35 36 341 286 362 FA_X1 $T=60660 45800 0 0 $X=60545 $Y=45685
X1636 178 298 324 325 35 36 122 360 362 FA_X1 $T=60850 48600 1 0 $X=60735 $Y=47085
X1637 203 30 219 341 35 36 123 360 362 FA_X1 $T=67500 48600 0 180 $X=64345 $Y=47085
X1638 92 299 326 354 35 36 125 285 361 FA_X1 $T=65220 51400 1 0 $X=65105 $Y=49885
X1639 124 358 309 342 35 36 94 360 362 FA_X1 $T=67500 48600 1 0 $X=67385 $Y=47085
X1640 181 300 132 350 35 36 359 360 361 FA_X1 $T=68640 48600 0 0 $X=68525 $Y=48485
X1641 183 359 214 151 35 36 126 360 361 FA_X1 $T=71680 48600 0 0 $X=71565 $Y=48485
X1642 96 343 133 153 35 36 344 360 362 FA_X1 $T=74910 48600 1 0 $X=74795 $Y=47085
X1643 186 215 185 152 35 36 343 286 362 FA_X1 $T=78330 45800 1 180 $X=75175 $Y=45685
X1644 300 32 220 211 35 36 327 285 361 FA_X1 $T=77190 51400 1 0 $X=77075 $Y=49885
X1645 97 356 189 105 35 36 301 286 362 FA_X1 $T=78330 45800 0 0 $X=78215 $Y=45685
X1646 127 301 344 212 35 36 187 360 361 FA_X1 $T=81750 48600 1 180 $X=78595 $Y=48485
X1647 188 33 327 155 35 36 345 285 361 FA_X1 $T=80230 51400 1 0 $X=80115 $Y=49885
X1648 98 302 328 355 35 36 101 360 362 FA_X1 $T=81750 48600 1 0 $X=81635 $Y=47085
X1649 99 345 190 158 35 36 356 360 361 FA_X1 $T=81750 48600 0 0 $X=81635 $Y=48485
X1650 351 69 36 290 11 165 35 286 362 OAI22_X1 $T=23230 45800 1 180 $X=22165 $Y=45685
X1651 139 35 106 66 36 315 360 361 NOR3_X1 $T=20950 48600 1 180 $X=20075 $Y=48485
X1652 25 35 85 147 36 82 360 361 NOR3_X1 $T=54770 48600 1 180 $X=53895 $Y=48485
X1654 37 35 289 63 135 304 36 285 361 NOR4_X1 $T=10500 51400 0 180 $X=9435 $Y=49885
X1655 38 35 64 159 161 160 36 286 362 NOR4_X1 $T=12400 45800 0 0 $X=12285 $Y=45685
X1656 136 35 9 163 62 162 36 360 361 NOR4_X1 $T=14680 48600 1 180 $X=13615 $Y=48485
X1657 143 35 167 168 169 316 36 286 362 NOR4_X1 $T=32160 45800 0 0 $X=32045 $Y=45685
X1658 289 48 36 35 360 361 INV_X2 $T=10690 48600 0 0 $X=10575 $Y=48485
X1659 63 77 36 35 285 361 INV_X2 $T=11070 51400 1 0 $X=10955 $Y=49885
X1660 9 164 36 35 360 362 INV_X2 $T=15060 48600 1 0 $X=14945 $Y=47085
X1661 144 49 36 35 286 362 INV_X2 $T=43940 45800 0 0 $X=43825 $Y=45685
X1662 12 14 15 36 35 104 360 362 OR3_X1 $T=23990 48600 1 0 $X=23875 $Y=47085
X1663 304 107 108 109 36 35 314 360 361 AND4_X1 $T=12590 48600 0 0 $X=12475 $Y=48485
.ENDS
***************************************
.SUBCKT ICV_14 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 30 31 32 33 34 35 36 37 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122
+ 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142
+ 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162
+ 163 164 165 166 167 168 169 170 171 172 173 227 228
** N=307 EP=173 IP=2790 FDC=1504
X919 271 4 26 25 97 305 306 DFF_X1 $T=1000 43000 1 0 $X=885 $Y=41485
X920 5 4 26 25 98 305 307 DFF_X1 $T=1760 43000 0 0 $X=1645 $Y=42885
X921 272 6 26 25 27 228 307 DFF_X1 $T=2900 45800 1 0 $X=2785 $Y=44285
X922 273 4 26 25 32 305 306 DFF_X1 $T=4230 43000 1 0 $X=4115 $Y=41485
X923 274 6 26 25 41 227 306 DFF_X1 $T=21140 40200 0 0 $X=21025 $Y=40085
X924 231 6 26 25 257 305 307 DFF_X1 $T=22470 43000 0 0 $X=22355 $Y=42885
X925 19 6 26 25 46 228 307 DFF_X1 $T=39380 45800 1 0 $X=39265 $Y=44285
X926 99 6 26 25 72 305 307 DFF_X1 $T=41090 43000 0 0 $X=40975 $Y=42885
X927 20 6 26 25 73 227 306 DFF_X1 $T=42420 40200 0 0 $X=42305 $Y=40085
X928 21 6 26 25 100 305 306 DFF_X1 $T=42610 43000 1 0 $X=42495 $Y=41485
X1049 250 26 25 272 228 307 CLKBUF_X1 $T=1000 45800 1 0 $X=885 $Y=44285
X1050 287 26 25 271 228 307 CLKBUF_X1 $T=1570 45800 1 0 $X=1455 $Y=44285
X1051 251 26 25 101 305 307 CLKBUF_X1 $T=6510 43000 0 0 $X=6395 $Y=42885
X1052 252 26 25 274 227 306 CLKBUF_X1 $T=8790 40200 0 0 $X=8675 $Y=40085
X1053 288 26 25 231 305 307 CLKBUF_X1 $T=9930 43000 0 0 $X=9815 $Y=42885
X1344 64 1 26 25 287 305 307 AND2_X1 $T=1000 43000 0 0 $X=885 $Y=42885
X1345 64 3 26 25 273 227 306 AND2_X1 $T=2900 40200 1 180 $X=2025 $Y=40085
X1346 28 2 26 25 250 228 307 AND2_X1 $T=2140 45800 1 0 $X=2025 $Y=44285
X1347 28 7 26 25 251 305 307 AND2_X1 $T=7840 43000 1 180 $X=6965 $Y=42885
X1348 28 8 26 25 288 305 307 AND2_X1 $T=9170 43000 0 0 $X=9055 $Y=42885
X1349 28 9 26 25 252 227 306 AND2_X1 $T=10120 40200 1 180 $X=9245 $Y=40085
X1350 64 11 26 25 129 228 307 AND2_X1 $T=9930 45800 1 0 $X=9815 $Y=44285
X1365 17 26 25 68 228 307 INV_X1 $T=22090 45800 1 0 $X=21975 $Y=44285
X1366 117 26 25 74 305 306 INV_X1 $T=48500 43000 1 0 $X=48385 $Y=41485
X1367 72 26 25 52 305 307 INV_X1 $T=49450 43000 0 0 $X=49335 $Y=42885
X1368 46 26 25 85 228 307 INV_X1 $T=51160 45800 1 0 $X=51045 $Y=44285
X1479 77 25 49 245 26 305 307 NOR2_X1 $T=13160 43000 0 0 $X=13045 $Y=42885
X1480 78 25 33 254 26 305 307 NOR2_X1 $T=14680 43000 0 0 $X=14565 $Y=42885
X1481 22 25 66 229 26 305 306 NOR2_X1 $T=16770 43000 1 0 $X=16655 $Y=41485
X1482 42 25 56 276 26 305 307 NOR2_X1 $T=20190 43000 1 180 $X=19505 $Y=42885
X1483 76 25 84 256 26 305 307 NOR2_X1 $T=20760 43000 1 180 $X=20075 $Y=42885
X1484 15 25 16 39 26 228 307 NOR2_X1 $T=22470 45800 1 0 $X=22355 $Y=44285
X1485 40 25 18 159 26 228 307 NOR2_X1 $T=24180 45800 1 0 $X=24065 $Y=44285
X1486 22 25 47 294 26 305 307 NOR2_X1 $T=30260 43000 1 180 $X=29575 $Y=42885
X1487 42 25 69 258 26 228 307 NOR2_X1 $T=30830 45800 0 180 $X=30145 $Y=44285
X1488 76 25 119 289 26 305 307 NOR2_X1 $T=31780 43000 1 180 $X=31095 $Y=42885
X1489 70 25 49 232 26 305 306 NOR2_X1 $T=33680 43000 1 0 $X=33565 $Y=41485
X1490 48 25 33 295 26 227 306 NOR2_X1 $T=36340 40200 0 0 $X=36225 $Y=40085
X1491 70 25 33 259 26 227 306 NOR2_X1 $T=40140 40200 0 0 $X=40025 $Y=40085
X1492 58 25 49 140 26 228 307 NOR2_X1 $T=45650 45800 1 0 $X=45535 $Y=44285
X1493 110 25 33 141 26 228 307 NOR2_X1 $T=47740 45800 0 180 $X=47055 $Y=44285
X1494 110 25 49 142 26 228 307 NOR2_X1 $T=48880 45800 1 0 $X=48765 $Y=44285
X1495 75 25 33 111 26 228 307 NOR2_X1 $T=50590 45800 1 0 $X=50475 $Y=44285
X1496 53 25 91 297 26 227 306 NOR2_X1 $T=51350 40200 1 180 $X=50665 $Y=40085
X1497 76 25 74 261 26 305 306 NOR2_X1 $T=51350 43000 0 180 $X=50665 $Y=41485
X1498 77 25 54 304 26 305 306 NOR2_X1 $T=52490 43000 1 0 $X=52375 $Y=41485
X1499 78 25 95 290 26 305 306 NOR2_X1 $T=53820 43000 1 0 $X=53705 $Y=41485
X1500 79 25 33 112 26 228 307 NOR2_X1 $T=54770 45800 0 180 $X=54085 $Y=44285
X1501 22 25 74 96 26 305 307 NOR2_X1 $T=55340 43000 0 0 $X=55225 $Y=42885
X1502 143 25 119 233 26 227 306 NOR2_X1 $T=55720 40200 0 0 $X=55605 $Y=40085
X1503 79 25 49 144 26 228 307 NOR2_X1 $T=57240 45800 1 0 $X=57125 $Y=44285
X1504 80 25 122 234 26 305 306 NOR2_X1 $T=58760 43000 1 0 $X=58645 $Y=41485
X1505 85 25 33 145 26 228 307 NOR2_X1 $T=59710 45800 0 180 $X=59025 $Y=44285
X1506 82 25 47 300 26 228 307 NOR2_X1 $T=59710 45800 1 0 $X=59595 $Y=44285
X1507 123 25 69 280 26 305 306 NOR2_X1 $T=60660 43000 1 0 $X=60545 $Y=41485
X1508 52 25 33 83 26 305 307 NOR2_X1 $T=61990 43000 1 180 $X=61305 $Y=42885
X1509 79 25 84 148 26 228 307 NOR2_X1 $T=61610 45800 1 0 $X=61495 $Y=44285
X1510 52 25 49 249 26 305 307 NOR2_X1 $T=61990 43000 0 0 $X=61875 $Y=42885
X1511 85 25 49 149 26 228 307 NOR2_X1 $T=62180 45800 1 0 $X=62065 $Y=44285
X1512 79 25 56 236 26 305 307 NOR2_X1 $T=63510 43000 0 0 $X=63395 $Y=42885
X1513 85 25 84 286 26 305 307 NOR2_X1 $T=64840 43000 0 0 $X=64725 $Y=42885
X1514 58 25 67 269 26 305 307 NOR2_X1 $T=67120 43000 0 0 $X=67005 $Y=42885
X1515 110 25 153 301 26 227 306 NOR2_X1 $T=68830 40200 1 180 $X=68145 $Y=40085
X1516 75 25 66 291 26 227 306 NOR2_X1 $T=68830 40200 0 0 $X=68715 $Y=40085
X1517 87 25 88 302 26 305 306 NOR2_X1 $T=71110 43000 1 0 $X=70995 $Y=41485
X1518 48 25 89 265 26 305 306 NOR2_X1 $T=71680 43000 1 0 $X=71565 $Y=41485
X1519 70 25 125 266 26 305 306 NOR2_X1 $T=73770 43000 0 180 $X=73085 $Y=41485
X1520 42 25 74 292 26 305 307 NOR2_X1 $T=73390 43000 0 0 $X=73275 $Y=42885
X1521 126 25 127 282 26 305 306 NOR2_X1 $T=75670 43000 1 0 $X=75555 $Y=41485
X1522 90 25 128 268 26 305 306 NOR2_X1 $T=76240 43000 1 0 $X=76125 $Y=41485
X1523 143 25 63 242 26 227 306 NOR2_X1 $T=78520 40200 0 0 $X=78405 $Y=40085
X1524 30 25 91 244 26 228 307 NOR2_X1 $T=81180 45800 1 0 $X=81065 $Y=44285
X1525 53 25 157 303 26 305 307 NOR2_X1 $T=82890 43000 0 0 $X=82775 $Y=42885
X1526 158 25 122 293 26 305 307 NOR2_X1 $T=83460 43000 0 0 $X=83345 $Y=42885
X1527 15 26 16 17 25 228 307 NAND2_X1 $T=21520 45800 1 0 $X=21405 $Y=44285
X1528 40 26 18 133 25 228 307 NAND2_X1 $T=25320 45800 0 180 $X=24635 $Y=44285
X1529 40 18 160 159 26 25 228 307 AOI21_X1 $T=26080 45800 0 180 $X=25205 $Y=44285
X1532 10 12 130 31 25 26 253 227 306 FA_X1 $T=10120 40200 0 0 $X=10005 $Y=40085
X1533 34 115 253 14 25 26 230 305 306 FA_X1 $T=16200 43000 0 180 $X=13045 $Y=41485
X1534 131 245 254 116 25 26 255 228 307 FA_X1 $T=15440 45800 1 0 $X=15325 $Y=44285
X1535 35 229 276 256 25 26 275 305 307 FA_X1 $T=16580 43000 0 0 $X=16465 $Y=42885
X1536 36 230 167 246 25 26 102 227 306 FA_X1 $T=18100 40200 0 0 $X=17985 $Y=40085
X1537 132 255 275 161 25 26 246 228 307 FA_X1 $T=21520 45800 0 180 $X=18365 $Y=44285
X1538 93 248 168 44 25 26 247 305 307 FA_X1 $T=26650 43000 0 0 $X=26535 $Y=42885
X1539 105 172 247 173 25 26 45 227 306 FA_X1 $T=27220 40200 0 0 $X=27105 $Y=40085
X1540 137 294 258 289 25 26 106 228 307 FA_X1 $T=27220 45800 1 0 $X=27105 $Y=44285
X1541 248 169 278 71 25 26 108 305 307 FA_X1 $T=35960 43000 0 0 $X=35845 $Y=42885
X1542 94 232 295 257 25 26 107 305 306 FA_X1 $T=39570 43000 0 180 $X=36415 $Y=41485
X1543 109 170 259 139 25 26 278 305 306 FA_X1 $T=42610 43000 0 180 $X=39455 $Y=41485
X1544 296 163 297 120 25 26 51 227 306 FA_X1 $T=45650 40200 0 0 $X=45535 $Y=40085
X1545 267 261 304 290 25 26 299 305 307 FA_X1 $T=52300 43000 0 0 $X=52185 $Y=42885
X1546 298 299 165 164 25 26 113 227 306 FA_X1 $T=52680 40200 0 0 $X=52565 $Y=40085
X1547 55 262 279 296 25 26 235 305 306 FA_X1 $T=55720 43000 1 0 $X=55605 $Y=41485
X1548 262 233 23 121 25 26 81 227 306 FA_X1 $T=56290 40200 0 0 $X=56175 $Y=40085
X1549 279 234 300 280 25 26 146 305 307 FA_X1 $T=58380 43000 0 0 $X=58265 $Y=42885
X1550 240 235 147 124 25 26 263 227 306 FA_X1 $T=59330 40200 0 0 $X=59215 $Y=40085
X1551 86 263 151 284 25 26 57 227 306 FA_X1 $T=62370 40200 0 0 $X=62255 $Y=40085
X1552 237 236 286 249 25 26 281 305 306 FA_X1 $T=62750 43000 1 0 $X=62635 $Y=41485
X1553 150 237 264 162 25 26 152 228 307 FA_X1 $T=62750 45800 1 0 $X=62635 $Y=44285
X1554 264 269 301 291 25 26 238 305 306 FA_X1 $T=65790 43000 1 0 $X=65675 $Y=41485
X1555 171 24 281 238 25 26 154 228 307 FA_X1 $T=68830 45800 1 0 $X=68715 $Y=44285
X1556 241 302 266 265 25 26 59 227 306 FA_X1 $T=69400 40200 0 0 $X=69285 $Y=40085
X1557 155 239 267 292 25 26 60 228 307 FA_X1 $T=71870 45800 1 0 $X=71755 $Y=44285
X1558 156 240 298 270 25 26 61 227 306 FA_X1 $T=75480 40200 0 0 $X=75365 $Y=40085
X1559 62 241 283 166 25 26 114 228 307 FA_X1 $T=78140 45800 1 0 $X=78025 $Y=44285
X1560 283 242 268 282 25 26 243 305 306 FA_X1 $T=78710 43000 1 0 $X=78595 $Y=41485
X1561 270 243 92 285 25 26 284 305 306 FA_X1 $T=81750 43000 1 0 $X=81635 $Y=41485
X1562 239 244 303 293 25 26 285 228 307 FA_X1 $T=81750 45800 1 0 $X=81635 $Y=44285
X1563 46 25 41 257 26 138 228 307 NOR3_X1 $T=33300 45800 1 0 $X=33185 $Y=44285
X1570 117 25 13 32 97 65 26 305 307 NOR4_X1 $T=12210 43000 0 0 $X=12095 $Y=42885
X1571 118 25 43 134 135 277 26 305 307 NOR4_X1 $T=25700 43000 0 0 $X=25585 $Y=42885
X1572 72 25 100 73 139 260 26 305 307 NOR4_X1 $T=44320 43000 0 0 $X=44205 $Y=42885
X1574 31 153 26 25 305 307 INV_X2 $T=11070 43000 1 180 $X=10385 $Y=42885
X1575 116 30 26 25 228 307 INV_X2 $T=11260 45800 0 180 $X=10575 $Y=44285
X1576 37 67 26 25 305 307 INV_X2 $T=21900 43000 0 0 $X=21785 $Y=42885
X1577 97 47 26 25 227 306 INV_X2 $T=26650 40200 0 0 $X=26535 $Y=40085
X1578 257 58 26 25 305 307 INV_X2 $T=39000 43000 0 0 $X=38885 $Y=42885
X1579 41 110 26 25 228 307 INV_X2 $T=42610 45800 1 0 $X=42495 $Y=44285
X1580 73 75 26 25 305 307 INV_X2 $T=46410 43000 0 0 $X=46295 $Y=42885
X1581 13 95 26 25 305 307 INV_X2 $T=47550 43000 0 0 $X=47435 $Y=42885
X1582 50 54 26 25 305 306 INV_X2 $T=47930 43000 1 0 $X=47815 $Y=41485
X1583 100 79 26 25 305 307 INV_X2 $T=48120 43000 0 0 $X=48005 $Y=42885
X1584 103 104 277 260 26 25 136 228 307 AND4_X1 $T=26080 45800 1 0 $X=25965 $Y=44285
.ENDS
***************************************
.SUBCKT ICV_15
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 37 38 39 40 41
+ 42 43 44 45 46 47 48 49 50 51 52 53 54 55 57 58 59 60 61 62
+ 63 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82 83
+ 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102 103
+ 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121 122 123
+ 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141 142 143
+ 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161 162 163
+ 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181 182 183
+ 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201 202 203
+ 204 205 206 207 208 209 210 211 212 213 214 215 216 217 218 219 220 221 222 223
+ 224 225 226 227 251 252
** N=473 EP=226 IP=5106 FDC=3182
X1722 329 6 38 37 85 467 471 DFF_X1 $T=1000 31800 1 0 $X=885 $Y=30285
X1723 398 6 38 37 384 468 473 DFF_X1 $T=1000 34600 1 0 $X=885 $Y=33085
X1724 399 6 38 37 83 468 472 DFF_X1 $T=2520 34600 0 0 $X=2405 $Y=34485
X1725 254 6 38 37 134 251 470 DFF_X1 $T=3280 40200 1 0 $X=3165 $Y=38685
X1726 255 6 38 37 40 469 470 DFF_X1 $T=3470 37400 0 0 $X=3355 $Y=37285
X1727 383 6 38 37 86 252 471 DFF_X1 $T=4230 29000 0 0 $X=4115 $Y=28885
X1728 385 6 38 37 41 468 473 DFF_X1 $T=4230 34600 1 0 $X=4115 $Y=33085
X1729 400 6 38 37 135 469 470 DFF_X1 $T=16200 37400 0 0 $X=16085 $Y=37285
X1730 133 6 38 37 51 467 473 DFF_X1 $T=16960 31800 0 0 $X=16845 $Y=31685
X1731 14 6 38 37 92 468 472 DFF_X1 $T=17530 34600 0 0 $X=17415 $Y=34485
X1732 124 16 38 37 95 251 470 DFF_X1 $T=19240 40200 1 0 $X=19125 $Y=38685
X1988 302 38 37 383 469 472 CLKBUF_X1 $T=1760 37400 1 0 $X=1645 $Y=35885
X1989 303 38 37 399 469 470 CLKBUF_X1 $T=1760 37400 0 0 $X=1645 $Y=37285
X1990 330 38 37 254 251 470 CLKBUF_X1 $T=1950 40200 1 0 $X=1835 $Y=38685
X1991 428 38 37 398 469 472 CLKBUF_X1 $T=2900 37400 0 180 $X=2215 $Y=35885
X1992 253 38 37 255 469 472 CLKBUF_X1 $T=2900 37400 1 0 $X=2785 $Y=35885
X1993 304 38 37 385 469 472 CLKBUF_X1 $T=4230 37400 1 0 $X=4115 $Y=35885
X1994 402 38 37 400 469 472 CLKBUF_X1 $T=6320 37400 1 0 $X=6205 $Y=35885
X1995 431 38 37 141 251 470 CLKBUF_X1 $T=36720 40200 1 0 $X=36605 $Y=38685
X1996 273 38 37 174 251 470 CLKBUF_X1 $T=39950 40200 1 0 $X=39835 $Y=38685
X1997 382 38 37 175 469 470 CLKBUF_X1 $T=40520 37400 0 0 $X=40405 $Y=37285
X1998 346 38 37 176 469 470 CLKBUF_X1 $T=42230 37400 0 0 $X=42115 $Y=37285
X2426 39 3 38 37 82 468 472 AND2_X1 $T=1760 34600 1 180 $X=885 $Y=34485
X2427 39 1 38 37 302 469 472 AND2_X1 $T=1000 37400 1 0 $X=885 $Y=35885
X2428 39 2 38 37 303 469 470 AND2_X1 $T=1000 37400 0 0 $X=885 $Y=37285
X2429 39 4 38 37 329 251 470 AND2_X1 $T=1760 40200 0 180 $X=885 $Y=38685
X2430 39 5 38 37 428 468 472 AND2_X1 $T=1760 34600 0 0 $X=1645 $Y=34485
X2431 39 7 38 37 330 251 470 AND2_X1 $T=2520 40200 1 0 $X=2405 $Y=38685
X2432 39 8 38 37 253 469 470 AND2_X1 $T=2710 37400 0 0 $X=2595 $Y=37285
X2433 39 9 38 37 304 469 472 AND2_X1 $T=3470 37400 1 0 $X=3355 $Y=35885
X2434 39 10 38 37 402 469 472 AND2_X1 $T=6890 37400 1 0 $X=6775 $Y=35885
X2435 93 15 38 37 53 252 471 AND2_X1 $T=19620 29000 0 0 $X=19505 $Y=28885
X2436 69 19 38 37 431 251 470 AND2_X1 $T=37290 40200 1 0 $X=37175 $Y=38685
X2437 69 22 38 37 273 251 470 AND2_X1 $T=41280 40200 0 180 $X=40405 $Y=38685
X2438 69 24 38 37 382 469 470 AND2_X1 $T=41850 37400 1 180 $X=40975 $Y=37285
X2439 69 25 38 37 346 469 470 AND2_X1 $T=42800 37400 0 0 $X=42685 $Y=37285
X2440 189 28 38 37 30 252 471 AND2_X1 $T=52490 29000 1 180 $X=51615 $Y=28885
X2473 357 38 37 73 252 471 INV_X1 $T=55530 29000 1 180 $X=55035 $Y=28885
X2508 28 453 27 38 37 354 252 471 HA_X1 $T=51730 29000 1 180 $X=49715 $Y=28885
X2509 389 354 280 38 37 191 467 473 HA_X1 $T=53630 31800 0 0 $X=53515 $Y=31685
X2691 44 37 21 441 38 468 472 NOR2_X1 $T=10690 34600 1 180 $X=10005 $Y=34485
X2692 46 37 12 442 38 469 472 NOR2_X1 $T=11260 37400 0 180 $X=10575 $Y=35885
X2693 108 37 45 256 38 469 470 NOR2_X1 $T=11070 37400 0 0 $X=10955 $Y=37285
X2694 106 37 45 258 38 467 473 NOR2_X1 $T=11830 31800 0 0 $X=11715 $Y=31685
X2695 108 37 91 332 38 252 471 NOR2_X1 $T=13160 29000 1 180 $X=12475 $Y=28885
X2696 46 37 48 259 38 468 472 NOR2_X1 $T=12590 34600 0 0 $X=12475 $Y=34485
X2697 106 37 47 331 38 469 470 NOR2_X1 $T=13160 37400 1 180 $X=12475 $Y=37285
X2698 59 37 47 305 38 467 473 NOR2_X1 $T=13920 31800 1 180 $X=13235 $Y=31685
X2699 181 37 102 306 38 468 472 NOR2_X1 $T=14490 34600 1 180 $X=13805 $Y=34485
X2700 50 37 91 404 38 469 472 NOR2_X1 $T=16770 37400 0 180 $X=16085 $Y=35885
X2701 44 37 12 333 38 251 470 NOR2_X1 $T=18670 40200 1 0 $X=18555 $Y=38685
X2702 15 37 93 55 38 467 471 NOR2_X1 $T=20190 31800 0 180 $X=19505 $Y=30285
X2703 44 37 54 430 38 467 473 NOR2_X1 $T=23610 31800 1 180 $X=22925 $Y=31685
X2704 44 37 71 334 38 469 470 NOR2_X1 $T=24370 37400 0 0 $X=24255 $Y=37285
X2705 46 37 54 335 38 469 472 NOR2_X1 $T=25890 37400 0 180 $X=25205 $Y=35885
X2706 59 37 58 264 38 469 472 NOR2_X1 $T=27790 37400 0 180 $X=27105 $Y=35885
X2707 161 37 21 61 38 252 471 NOR2_X1 $T=28360 29000 0 0 $X=28245 $Y=28885
X2708 98 37 62 336 38 251 470 NOR2_X1 $T=29880 40200 1 0 $X=29765 $Y=38685
X2709 99 37 100 337 38 469 472 NOR2_X1 $T=30450 37400 1 0 $X=30335 $Y=35885
X2710 65 37 45 267 38 467 471 NOR2_X1 $T=34250 31800 0 180 $X=33565 $Y=30285
X2711 101 37 47 338 38 252 471 NOR2_X1 $T=35390 29000 1 180 $X=34705 $Y=28885
X2712 67 37 48 270 38 468 473 NOR2_X1 $T=35580 34600 1 0 $X=35465 $Y=33085
X2713 70 37 48 447 38 467 473 NOR2_X1 $T=37100 31800 1 180 $X=36415 $Y=31685
X2714 101 37 91 448 38 469 472 NOR2_X1 $T=36720 37400 1 0 $X=36605 $Y=35885
X2715 65 37 102 315 38 468 473 NOR2_X1 $T=37480 34600 1 0 $X=37365 $Y=33085
X2716 161 37 103 271 38 251 470 NOR2_X1 $T=38050 40200 1 0 $X=37935 $Y=38685
X2717 108 37 20 340 38 252 471 NOR2_X1 $T=39000 29000 1 180 $X=38315 $Y=28885
X2718 65 37 91 388 38 467 473 NOR2_X1 $T=38620 31800 0 0 $X=38505 $Y=31685
X2719 70 37 12 411 38 251 470 NOR2_X1 $T=39380 40200 0 180 $X=38695 $Y=38685
X2720 67 37 102 272 38 467 473 NOR2_X1 $T=39760 31800 1 180 $X=39075 $Y=31685
X2721 162 37 21 341 38 468 472 NOR2_X1 $T=39190 34600 0 0 $X=39075 $Y=34485
X2722 101 37 45 198 38 251 470 NOR2_X1 $T=39380 40200 1 0 $X=39265 $Y=38685
X2723 101 37 68 316 38 468 472 NOR2_X1 $T=39760 34600 0 0 $X=39645 $Y=34485
X2724 79 37 163 449 38 467 473 NOR2_X1 $T=41090 31800 0 0 $X=40975 $Y=31685
X2725 116 37 58 318 38 468 472 NOR2_X1 $T=41660 34600 0 0 $X=41545 $Y=34485
X2726 98 37 121 276 38 251 470 NOR2_X1 $T=44700 40200 1 0 $X=44585 $Y=38685
X2727 70 37 71 348 38 469 472 NOR2_X1 $T=44890 37400 1 0 $X=44775 $Y=35885
X2728 161 37 105 349 38 469 472 NOR2_X1 $T=46790 37400 0 180 $X=46105 $Y=35885
X2729 162 37 173 432 38 469 470 NOR2_X1 $T=47170 37400 1 180 $X=46485 $Y=37285
X2730 67 37 54 451 38 468 472 NOR2_X1 $T=47550 34600 1 180 $X=46865 $Y=34485
X2731 65 37 72 352 38 468 473 NOR2_X1 $T=47740 34600 0 180 $X=47055 $Y=33085
X2732 106 37 107 200 38 251 470 NOR2_X1 $T=47170 40200 1 0 $X=47055 $Y=38685
X2733 99 37 121 109 38 251 470 NOR2_X1 $T=49640 40200 0 180 $X=48955 $Y=38685
X2734 108 37 110 464 38 468 473 NOR2_X1 $T=49260 34600 1 0 $X=49145 $Y=33085
X2735 50 37 20 353 38 468 472 NOR2_X1 $T=49450 34600 0 0 $X=49335 $Y=34485
X2736 30 37 166 190 38 252 471 NOR2_X1 $T=54010 29000 0 0 $X=53895 $Y=28885
X2737 389 37 279 357 38 252 471 NOR2_X1 $T=56100 29000 1 180 $X=55415 $Y=28885
X2738 65 37 68 75 38 469 470 NOR2_X1 $T=57620 37400 0 0 $X=57505 $Y=37285
X2739 114 37 12 283 38 467 473 NOR2_X1 $T=58570 31800 0 0 $X=58455 $Y=31685
X2740 67 37 72 201 38 251 470 NOR2_X1 $T=59140 40200 0 180 $X=58455 $Y=38685
X2741 76 37 102 434 38 467 473 NOR2_X1 $T=59900 31800 0 0 $X=59785 $Y=31685
X2742 101 37 163 323 38 251 470 NOR2_X1 $T=60280 40200 1 0 $X=60165 $Y=38685
X2743 78 37 48 358 38 467 471 NOR2_X1 $T=61420 31800 0 180 $X=60735 $Y=30285
X2744 114 37 68 284 38 467 471 NOR2_X1 $T=61420 31800 1 0 $X=61305 $Y=30285
X2745 79 37 58 457 38 469 472 NOR2_X1 $T=62750 37400 0 180 $X=62065 $Y=35885
X2746 81 37 62 392 38 468 472 NOR2_X1 $T=62940 34600 1 180 $X=62255 $Y=34485
X2747 34 37 103 324 38 467 473 NOR2_X1 $T=63510 31800 1 180 $X=62825 $Y=31685
X2748 118 37 21 359 38 468 472 NOR2_X1 $T=63510 34600 1 180 $X=62825 $Y=34485
X2749 116 37 100 360 38 469 470 NOR2_X1 $T=63510 37400 1 180 $X=62825 $Y=37285
X2750 76 37 58 325 38 467 471 NOR2_X1 $T=63700 31800 0 180 $X=63015 $Y=30285
X2751 78 37 163 326 38 467 471 NOR2_X1 $T=63700 31800 1 0 $X=63585 $Y=30285
X2752 76 37 91 436 38 469 472 NOR2_X1 $T=64650 37400 1 0 $X=64535 $Y=35885
X2753 101 37 115 286 38 468 473 NOR2_X1 $T=64840 34600 1 0 $X=64725 $Y=33085
X2754 114 37 48 327 38 469 472 NOR2_X1 $T=65220 37400 1 0 $X=65105 $Y=35885
X2755 116 37 105 435 38 468 473 NOR2_X1 $T=66930 34600 0 180 $X=66245 $Y=33085
X2756 162 37 20 419 38 467 473 NOR2_X1 $T=67120 31800 1 180 $X=66435 $Y=31685
X2757 78 37 102 459 38 469 472 NOR2_X1 $T=67310 37400 0 180 $X=66625 $Y=35885
X2758 79 37 121 362 38 468 472 NOR2_X1 $T=68070 34600 1 180 $X=67385 $Y=34485
X2759 118 37 12 363 38 251 470 NOR2_X1 $T=68830 40200 0 180 $X=68145 $Y=38685
X2760 70 37 20 288 38 468 473 NOR2_X1 $T=69400 34600 1 0 $X=69285 $Y=33085
X2761 81 37 103 461 38 468 472 NOR2_X1 $T=69970 34600 1 180 $X=69285 $Y=34485
X2762 67 37 110 364 38 468 473 NOR2_X1 $T=70540 34600 0 180 $X=69855 $Y=33085
X2763 34 37 21 460 38 468 472 NOR2_X1 $T=69970 34600 0 0 $X=69855 $Y=34485
X2764 65 37 107 437 38 467 473 NOR2_X1 $T=72250 31800 1 180 $X=71565 $Y=31685
X2765 67 37 20 328 38 468 473 NOR2_X1 $T=72820 34600 1 0 $X=72705 $Y=33085
X2766 65 37 110 394 38 467 473 NOR2_X1 $T=73770 31800 0 0 $X=73655 $Y=31685
X2767 101 37 107 294 38 251 470 NOR2_X1 $T=73960 40200 1 0 $X=73845 $Y=38685
X2768 101 37 110 292 38 467 473 NOR2_X1 $T=74910 31800 1 180 $X=74225 $Y=31685
X2769 79 37 107 373 38 467 473 NOR2_X1 $T=75860 31800 0 0 $X=75745 $Y=31685
X2770 79 37 115 371 38 251 470 NOR2_X1 $T=75860 40200 1 0 $X=75745 $Y=38685
X2771 116 37 115 438 38 467 473 NOR2_X1 $T=77190 31800 0 0 $X=77075 $Y=31685
X2772 116 37 121 396 38 251 470 NOR2_X1 $T=77950 40200 1 0 $X=77835 $Y=38685
X2773 81 37 105 297 38 469 470 NOR2_X1 $T=79090 37400 0 0 $X=78975 $Y=37285
X2774 34 37 173 377 38 469 470 NOR2_X1 $T=79660 37400 0 0 $X=79545 $Y=37285
X2775 114 37 173 298 38 252 471 NOR2_X1 $T=81180 29000 1 180 $X=80495 $Y=28885
X2776 81 37 121 300 38 468 472 NOR2_X1 $T=80610 34600 0 0 $X=80495 $Y=34485
X2777 118 37 71 425 38 251 470 NOR2_X1 $T=82130 40200 0 180 $X=81445 $Y=38685
X2778 114 37 54 301 38 251 470 NOR2_X1 $T=82130 40200 1 0 $X=82015 $Y=38685
X2779 34 37 105 379 38 469 472 NOR2_X1 $T=82510 37400 1 0 $X=82395 $Y=35885
X2780 76 37 54 426 38 467 471 NOR2_X1 $T=83460 31800 1 0 $X=83345 $Y=30285
X2781 78 37 71 462 38 467 473 NOR2_X1 $T=84030 31800 1 180 $X=83345 $Y=31685
X2782 76 37 68 380 38 251 470 NOR2_X1 $T=83460 40200 1 0 $X=83345 $Y=38685
X2783 78 37 72 381 38 251 470 NOR2_X1 $T=84600 40200 0 180 $X=83915 $Y=38685
X2784 78 37 54 427 38 252 471 NOR2_X1 $T=84790 29000 1 180 $X=84105 $Y=28885
X2785 118 37 173 440 38 468 472 NOR2_X1 $T=84790 34600 1 180 $X=84105 $Y=34485
X2786 38 390 454 32 37 252 471 XNOR2_X1 $T=56860 29000 0 0 $X=56745 $Y=28885
X2787 169 38 455 147 37 252 471 NAND2_X1 $T=58950 29000 0 0 $X=58835 $Y=28885
X2788 389 279 390 357 38 37 252 471 AOI21_X1 $T=56860 29000 1 180 $X=55985 $Y=28885
X2800 389 279 37 125 30 38 73 112 252 471 AOI221_X1 $T=54010 29000 1 180 $X=52755 $Y=28885
X2801 136 215 386 429 37 38 401 467 471 FA_X1 $T=9930 31800 0 180 $X=6775 $Y=30285
X2802 429 11 177 332 37 38 257 252 471 FA_X1 $T=7460 29000 0 0 $X=7345 $Y=28885
X2803 260 42 441 442 37 38 403 469 472 FA_X1 $T=7650 37400 1 0 $X=7535 $Y=35885
X2804 43 256 331 87 37 38 261 251 470 FA_X1 $T=9170 40200 1 0 $X=9055 $Y=38685
X2805 443 257 403 202 37 38 88 467 471 FA_X1 $T=9930 31800 1 0 $X=9815 $Y=30285
X2806 386 258 305 178 37 38 89 468 473 FA_X1 $T=10690 34600 1 0 $X=10575 $Y=33085
X2807 126 259 306 404 37 38 307 469 472 FA_X1 $T=11260 37400 1 0 $X=11145 $Y=35885
X2808 196 260 157 333 37 38 308 251 470 FA_X1 $T=12210 40200 1 0 $X=12095 $Y=38685
X2809 179 216 212 211 37 38 183 467 471 FA_X1 $T=12970 31800 1 0 $X=12855 $Y=30285
X2810 180 261 307 308 37 38 262 469 470 FA_X1 $T=13160 37400 0 0 $X=13045 $Y=37285
X2811 90 203 443 401 37 38 405 467 473 FA_X1 $T=13920 31800 0 0 $X=13805 $Y=31685
X2812 182 13 405 262 37 38 52 468 472 FA_X1 $T=14490 34600 0 0 $X=14375 $Y=34485
X2813 138 444 384 430 37 38 407 467 471 FA_X1 $T=21140 31800 1 0 $X=21025 $Y=30285
X2814 444 17 334 335 37 38 184 469 472 FA_X1 $T=22280 37400 1 0 $X=22165 $Y=35885
X2815 309 263 96 204 37 38 406 251 470 FA_X1 $T=25510 40200 0 180 $X=22355 $Y=38685
X2816 197 205 310 227 37 38 139 468 473 FA_X1 $T=23420 34600 1 0 $X=23305 $Y=33085
X2817 263 264 337 336 37 38 408 469 470 FA_X1 $T=24940 37400 0 0 $X=24825 $Y=37285
X2818 57 206 407 309 37 38 266 252 471 FA_X1 $T=25320 29000 0 0 $X=25205 $Y=28885
X2819 310 217 265 311 37 38 97 468 472 FA_X1 $T=26270 34600 0 0 $X=26155 $Y=34485
X2820 127 207 387 160 37 38 265 467 471 FA_X1 $T=27600 31800 1 0 $X=27485 $Y=30285
X2821 311 266 208 312 37 38 140 468 472 FA_X1 $T=29310 34600 0 0 $X=29195 $Y=34485
X2822 387 213 445 409 37 38 60 467 473 FA_X1 $T=29880 31800 0 0 $X=29765 $Y=31685
X2823 226 267 338 95 37 38 409 467 471 FA_X1 $T=33680 31800 0 180 $X=30525 $Y=30285
X2824 314 269 342 408 37 38 63 469 470 FA_X1 $T=36340 37400 1 180 $X=33185 $Y=37285
X2825 128 268 218 344 37 38 445 467 473 FA_X1 $T=33490 31800 0 0 $X=33375 $Y=31685
X2826 268 18 313 339 37 38 446 469 472 FA_X1 $T=33680 37400 1 0 $X=33565 $Y=35885
X2827 312 314 406 446 37 38 185 251 470 FA_X1 $T=33680 40200 1 0 $X=33565 $Y=38685
X2828 410 219 186 340 37 38 142 252 471 FA_X1 $T=35390 29000 0 0 $X=35275 $Y=28885
X2829 313 270 315 448 37 38 269 468 472 FA_X1 $T=36150 34600 0 0 $X=36035 $Y=34485
X2830 339 271 341 411 37 38 342 469 472 FA_X1 $T=37290 37400 1 0 $X=37175 $Y=35885
X2831 344 447 272 388 37 38 66 467 471 FA_X1 $T=41850 31800 0 180 $X=38695 $Y=30285
X2832 274 316 449 318 37 38 275 468 473 FA_X1 $T=39570 34600 1 0 $X=39455 $Y=33085
X2833 199 274 345 450 37 38 320 469 472 FA_X1 $T=40330 37400 1 0 $X=40215 $Y=35885
X2834 343 23 187 164 37 38 143 252 471 FA_X1 $T=40710 29000 0 0 $X=40595 $Y=28885
X2835 317 220 319 320 37 38 277 467 471 FA_X1 $T=41850 31800 1 0 $X=41735 $Y=30285
X2836 319 275 350 412 37 38 144 467 473 FA_X1 $T=43560 31800 0 0 $X=43445 $Y=31685
X2837 450 276 349 432 37 38 412 469 470 FA_X1 $T=43560 37400 0 0 $X=43445 $Y=37285
X2838 463 466 221 209 37 38 278 252 471 FA_X1 $T=43750 29000 0 0 $X=43635 $Y=28885
X2839 345 348 451 352 37 38 350 468 472 FA_X1 $T=43940 34600 0 0 $X=43825 $Y=34485
X2840 321 278 104 277 37 38 347 467 471 FA_X1 $T=47930 31800 0 180 $X=44775 $Y=30285
X2841 188 26 222 165 37 38 413 252 471 FA_X1 $T=46790 29000 0 0 $X=46675 $Y=28885
X2842 351 214 452 410 37 38 322 469 470 FA_X1 $T=47170 37400 0 0 $X=47055 $Y=37285
X2843 356 158 322 433 37 38 414 468 473 FA_X1 $T=49830 34600 1 0 $X=49715 $Y=33085
X2844 29 343 353 464 37 38 452 469 472 FA_X1 $T=53060 37400 0 180 $X=49905 $Y=35885
X2845 280 347 159 414 37 38 453 467 473 FA_X1 $T=50590 31800 0 0 $X=50475 $Y=31685
X2846 111 415 356 463 37 38 281 468 473 FA_X1 $T=52870 34600 1 0 $X=52755 $Y=33085
X2847 192 369 355 317 37 38 415 469 472 FA_X1 $T=56100 37400 0 180 $X=52945 $Y=35885
X2848 74 31 351 465 37 38 145 469 470 FA_X1 $T=54580 37400 0 0 $X=54465 $Y=37285
X2849 355 413 416 417 37 38 466 467 473 FA_X1 $T=55530 31800 0 0 $X=55415 $Y=31685
X2850 113 281 223 321 37 38 279 468 473 FA_X1 $T=55910 34600 1 0 $X=55795 $Y=33085
X2851 465 282 224 168 37 38 433 469 472 FA_X1 $T=56100 37400 1 0 $X=55985 $Y=35885
X2852 285 283 358 434 37 38 416 467 471 FA_X1 $T=57810 31800 1 0 $X=57695 $Y=30285
X2853 287 285 456 391 37 38 146 468 472 FA_X1 $T=61800 34600 1 180 $X=58645 $Y=34485
X2854 456 392 324 359 37 38 417 468 473 FA_X1 $T=58950 34600 1 0 $X=58835 $Y=33085
X2855 129 284 326 325 37 38 148 252 471 FA_X1 $T=59520 29000 0 0 $X=59405 $Y=28885
X2856 391 323 457 360 37 38 282 469 470 FA_X1 $T=59900 37400 0 0 $X=59785 $Y=37285
X2857 130 393 458 419 37 38 150 467 473 FA_X1 $T=63510 31800 0 0 $X=63395 $Y=31685
X2858 393 286 362 435 37 38 291 468 472 FA_X1 $T=63510 34600 0 0 $X=63395 $Y=34485
X2859 361 327 459 436 37 38 289 469 470 FA_X1 $T=63510 37400 0 0 $X=63395 $Y=37285
X2860 149 287 361 418 37 38 117 251 470 FA_X1 $T=65220 40200 1 0 $X=65105 $Y=38685
X2861 418 461 460 363 37 38 368 469 470 FA_X1 $T=66550 37400 0 0 $X=66435 $Y=37285
X2862 77 420 365 210 37 38 151 252 471 FA_X1 $T=68070 29000 0 0 $X=67955 $Y=28885
X2863 458 288 364 437 37 38 367 467 473 FA_X1 $T=68640 31800 0 0 $X=68525 $Y=31685
X2864 80 289 368 170 37 38 369 251 470 FA_X1 $T=70920 40200 1 0 $X=70805 $Y=38685
X2865 365 33 195 171 37 38 152 252 471 FA_X1 $T=71110 29000 0 0 $X=70995 $Y=28885
X2866 153 291 367 366 37 38 119 467 471 FA_X1 $T=74340 31800 0 180 $X=71185 $Y=30285
X2867 366 290 328 394 37 38 421 468 472 FA_X1 $T=71490 34600 0 0 $X=71375 $Y=34485
X2868 420 397 375 395 37 38 370 469 472 FA_X1 $T=73200 37400 1 0 $X=73085 $Y=35885
X2869 131 293 372 370 37 38 120 467 471 FA_X1 $T=77380 31800 0 180 $X=74225 $Y=30285
X2870 290 292 373 438 37 38 422 468 473 FA_X1 $T=75100 34600 1 0 $X=74985 $Y=33085
X2871 395 294 371 396 37 38 374 469 470 FA_X1 $T=76050 37400 0 0 $X=75935 $Y=37285
X2872 372 295 374 421 37 38 122 469 472 FA_X1 $T=76240 37400 1 0 $X=76125 $Y=35885
X2873 293 296 423 439 37 38 154 467 471 FA_X1 $T=77380 31800 1 0 $X=77265 $Y=30285
X2874 132 225 424 378 37 38 423 252 471 FA_X1 $T=77570 29000 0 0 $X=77455 $Y=28885
X2875 375 297 377 425 37 38 295 251 470 FA_X1 $T=78520 40200 1 0 $X=78405 $Y=38685
X2876 376 298 462 426 37 38 123 467 471 FA_X1 $T=80420 31800 1 0 $X=80305 $Y=30285
X2877 296 299 422 376 37 38 155 467 473 FA_X1 $T=80420 31800 0 0 $X=80305 $Y=31685
X2878 424 35 427 172 37 38 156 252 471 FA_X1 $T=81180 29000 0 0 $X=81065 $Y=28885
X2879 378 300 379 440 37 38 299 468 472 FA_X1 $T=81180 34600 0 0 $X=81065 $Y=34485
X2880 397 301 381 380 37 38 439 469 470 FA_X1 $T=81750 37400 0 0 $X=81635 $Y=37285
X2889 384 37 86 85 84 49 38 467 471 NOR4_X1 $T=6890 31800 0 180 $X=5825 $Y=30285
X2890 41 37 83 92 51 137 38 468 473 NOR4_X1 $T=16010 34600 1 0 $X=15895 $Y=33085
X2891 167 37 193 454 194 455 38 252 471 NOR4_X1 $T=58000 29000 0 0 $X=57885 $Y=28885
X2895 87 59 38 37 251 470 INV_X2 $T=9170 40200 0 180 $X=8485 $Y=38685
X2896 42 103 38 37 469 470 INV_X2 $T=9170 37400 0 0 $X=9055 $Y=37285
X2897 178 99 38 37 469 470 INV_X2 $T=9740 37400 0 0 $X=9625 $Y=37285
X2898 51 62 38 37 252 471 INV_X2 $T=19050 29000 0 0 $X=18935 $Y=28885
X2899 94 98 38 37 469 472 INV_X2 $T=20950 37400 1 0 $X=20835 $Y=35885
X2900 41 54 38 37 252 471 INV_X2 $T=22280 29000 0 0 $X=22165 $Y=28885
X2901 384 71 38 37 467 473 INV_X2 $T=24560 31800 0 0 $X=24445 $Y=31685
X2902 95 79 38 37 467 473 INV_X2 $T=32920 31800 0 0 $X=32805 $Y=31685
.ENDS
***************************************
.SUBCKT ICV_17 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 58 59 60 61
+ 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81
+ 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101
+ 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120 121
+ 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140 141
+ 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160 161
+ 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180 181
+ 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200 201
+ 202 203 204 205 206 207 208 209 210 211 212 213 214 215 240 241
** N=448 EP=216 IP=4791 FDC=2626
M0 19 303 31 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=4.3575e-14 PD=1.11e-06 PS=1.04e-06 $X=59705 $Y=22895 $D=1
M1 31 268 19 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=59895 $Y=22895 $D=1
M2 19 302 31 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=60085 $Y=22895 $D=1
M3 31 301 19 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=60275 $Y=22895 $D=1
M4 19 301 31 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=60465 $Y=22895 $D=1
M5 31 302 19 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=60655 $Y=22895 $D=1
M6 19 268 31 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=5.81e-14 AS=5.81e-14 PD=1.11e-06 PS=1.11e-06 $X=60845 $Y=22895 $D=1
M7 31 303 19 443 NMOS_VTL L=5e-08 W=4.15e-07 AD=4.3575e-14 AS=5.81e-14 PD=1.04e-06 PS=1.11e-06 $X=61035 $Y=22895 $D=1
M8 437 303 32 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=6.615e-14 PD=1.54e-06 PS=1.47e-06 $X=59705 $Y=22090 $D=0
M9 438 268 437 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=59895 $Y=22090 $D=0
M10 439 302 438 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=60085 $Y=22090 $D=0
M11 19 301 439 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=60275 $Y=22090 $D=0
M12 440 301 19 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=60465 $Y=22090 $D=0
M13 441 302 440 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=60655 $Y=22090 $D=0
M14 442 268 441 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=8.82e-14 AS=8.82e-14 PD=1.54e-06 PS=1.54e-06 $X=60845 $Y=22090 $D=0
M15 32 303 442 446 PMOS_VTL L=5e-08 W=6.3e-07 AD=6.615e-14 AS=8.82e-14 PD=1.47e-06 PS=1.54e-06 $X=61035 $Y=22090 $D=0
X1628 125 2 31 32 72 240 448 DFF_X1 $T=1000 29000 1 0 $X=885 $Y=27485
X2115 339 261 31 32 134 444 448 OR2_X1 $T=54200 26200 0 0 $X=54085 $Y=26085
X2299 96 20 31 32 301 445 241 AND2_X1 $T=54770 20600 0 180 $X=53895 $Y=19085
X2300 355 279 31 32 109 445 241 AND2_X1 $T=72060 20600 0 180 $X=71185 $Y=19085
X2325 336 18 372 260 31 32 443 446 OAI21_X1 $T=54770 23400 0 180 $X=53895 $Y=21885
X2326 340 262 393 338 31 32 444 447 OAI21_X1 $T=55150 26200 0 180 $X=54275 $Y=24685
X2327 344 21 166 341 31 32 240 448 OAI21_X1 $T=56480 29000 0 180 $X=55605 $Y=27485
X2328 68 274 406 269 31 32 445 446 OAI21_X1 $T=69400 20600 1 180 $X=68525 $Y=20485
X2329 113 30 124 27 31 32 445 241 OAI21_X1 $T=81940 20600 1 0 $X=81825 $Y=19085
X2330 411 31 32 262 443 447 INV_X1 $T=53440 23400 0 0 $X=53325 $Y=23285
X2331 63 31 32 341 240 448 INV_X1 $T=53630 29000 1 0 $X=53515 $Y=27485
X2332 337 31 32 338 444 447 INV_X1 $T=54010 26200 1 0 $X=53895 $Y=24685
X2333 393 31 32 344 444 448 INV_X1 $T=56480 26200 1 180 $X=55985 $Y=26085
X2334 414 31 32 343 445 446 INV_X1 $T=57240 20600 0 0 $X=57125 $Y=20485
X2335 100 31 32 415 445 241 INV_X1 $T=62750 20600 1 0 $X=62635 $Y=19085
X2336 428 31 32 121 445 241 INV_X1 $T=73580 20600 1 0 $X=73465 $Y=19085
X2369 332 330 16 31 32 95 443 446 HA_X1 $T=51540 23400 0 180 $X=49525 $Y=21885
X2370 336 93 17 31 32 335 445 241 HA_X1 $T=50590 20600 1 0 $X=50475 $Y=19085
X2371 347 186 273 31 32 67 445 241 HA_X1 $T=64650 20600 1 0 $X=64535 $Y=19085
X2372 279 360 280 31 32 122 445 446 HA_X1 $T=72250 20600 0 0 $X=72135 $Y=20485
X2373 110 361 281 31 32 360 445 446 HA_X1 $T=75860 20600 0 0 $X=75745 $Y=20485
X2374 417 436 29 31 32 281 445 446 HA_X1 $T=79850 20600 0 0 $X=79735 $Y=20485
X2547 74 32 88 418 31 445 446 NOR2_X1 $T=6130 20600 1 180 $X=5445 $Y=20485
X2548 83 32 4 306 31 445 446 NOR2_X1 $T=6890 20600 0 0 $X=6775 $Y=20485
X2549 74 32 4 407 31 443 446 NOR2_X1 $T=7080 23400 1 0 $X=6965 $Y=21885
X2550 75 32 37 36 31 240 448 NOR2_X1 $T=8980 29000 1 0 $X=8865 $Y=27485
X2551 82 32 35 286 31 443 447 NOR2_X1 $T=10500 23400 1 180 $X=9815 $Y=23285
X2552 80 32 37 243 31 445 446 NOR2_X1 $T=10690 20600 1 180 $X=10005 $Y=20485
X2553 49 32 79 77 31 240 448 NOR2_X1 $T=11830 29000 0 180 $X=11145 $Y=27485
X2554 38 32 46 420 31 443 447 NOR2_X1 $T=11830 23400 0 0 $X=11715 $Y=23285
X2555 52 32 79 307 31 445 446 NOR2_X1 $T=12020 20600 0 0 $X=11905 $Y=20485
X2556 12 32 8 310 31 443 446 NOR2_X1 $T=13160 23400 0 180 $X=12475 $Y=21885
X2557 74 32 142 246 31 443 446 NOR2_X1 $T=14300 23400 1 0 $X=14185 $Y=21885
X2558 49 32 37 367 31 445 241 NOR2_X1 $T=14870 20600 1 0 $X=14755 $Y=19085
X2559 80 32 79 421 31 445 241 NOR2_X1 $T=16010 20600 0 180 $X=15325 $Y=19085
X2560 52 32 8 404 31 445 446 NOR2_X1 $T=18100 20600 0 0 $X=17985 $Y=20485
X2561 12 32 35 314 31 444 448 NOR2_X1 $T=18670 26200 1 180 $X=17985 $Y=26085
X2562 75 32 10 289 31 443 447 NOR2_X1 $T=18860 23400 1 180 $X=18175 $Y=23285
X2563 83 32 146 313 31 443 447 NOR2_X1 $T=20380 23400 1 180 $X=19695 $Y=23285
X2564 82 32 46 384 31 444 447 NOR2_X1 $T=20000 26200 1 0 $X=19885 $Y=24685
X2565 83 32 22 385 31 444 447 NOR2_X1 $T=20570 26200 1 0 $X=20455 $Y=24685
X2566 75 32 13 290 31 444 448 NOR2_X1 $T=22470 26200 0 0 $X=22355 $Y=26085
X2567 49 32 85 316 31 240 448 NOR2_X1 $T=22850 29000 1 0 $X=22735 $Y=27485
X2568 38 32 142 248 31 240 448 NOR2_X1 $T=25700 29000 1 0 $X=25585 $Y=27485
X2569 66 32 10 319 31 444 448 NOR2_X1 $T=28740 26200 0 0 $X=28625 $Y=26085
X2570 75 32 22 432 31 444 447 NOR2_X1 $T=31970 26200 1 0 $X=31855 $Y=24685
X2571 52 32 117 253 31 445 446 NOR2_X1 $T=32540 20600 0 0 $X=32425 $Y=20485
X2572 82 32 4 409 31 445 446 NOR2_X1 $T=33110 20600 0 0 $X=32995 $Y=20485
X2573 50 32 46 87 31 445 241 NOR2_X1 $T=34060 20600 0 180 $X=33375 $Y=19085
X2574 12 32 88 433 31 443 446 NOR2_X1 $T=33490 23400 1 0 $X=33375 $Y=21885
X2575 80 32 85 321 31 240 448 NOR2_X1 $T=33870 29000 1 0 $X=33755 $Y=27485
X2576 49 32 13 434 31 444 447 NOR2_X1 $T=34060 26200 1 0 $X=33945 $Y=24685
X2577 89 32 65 390 31 443 446 NOR2_X1 $T=34820 23400 1 0 $X=34705 $Y=21885
X2578 103 32 13 322 31 445 446 NOR2_X1 $T=35010 20600 0 0 $X=34895 $Y=20485
X2579 102 32 22 368 31 445 446 NOR2_X1 $T=35580 20600 0 0 $X=35465 $Y=20485
X2580 115 32 105 255 31 443 447 NOR2_X1 $T=36150 23400 0 0 $X=36035 $Y=23285
X2581 50 32 99 292 31 443 447 NOR2_X1 $T=39000 23400 1 180 $X=38315 $Y=23285
X2582 52 32 54 53 31 240 448 NOR2_X1 $T=40710 29000 1 0 $X=40595 $Y=27485
X2583 60 32 117 295 31 444 448 NOR2_X1 $T=41470 26200 1 180 $X=40785 $Y=26085
X2584 12 32 55 161 31 444 448 NOR2_X1 $T=41470 26200 0 0 $X=41355 $Y=26085
X2585 91 32 88 326 31 444 447 NOR2_X1 $T=43750 26200 0 180 $X=43065 $Y=24685
X2586 82 32 145 56 31 444 448 NOR2_X1 $T=43940 26200 1 180 $X=43255 $Y=26085
X2587 62 32 4 369 31 444 448 NOR2_X1 $T=43940 26200 0 0 $X=43825 $Y=26085
X2588 92 32 142 257 31 445 446 NOR2_X1 $T=46410 20600 0 0 $X=46295 $Y=20485
X2589 26 32 146 328 31 445 446 NOR2_X1 $T=47930 20600 0 0 $X=47815 $Y=20485
X2590 94 32 10 370 31 445 446 NOR2_X1 $T=49070 20600 1 180 $X=48385 $Y=20485
X2591 92 32 146 259 31 443 446 NOR2_X1 $T=49640 23400 0 180 $X=48955 $Y=21885
X2592 60 32 88 258 31 240 448 NOR2_X1 $T=49450 29000 1 0 $X=49335 $Y=27485
X2593 26 32 10 299 31 444 447 NOR2_X1 $T=51540 26200 0 180 $X=50855 $Y=24685
X2594 91 32 4 300 31 240 448 NOR2_X1 $T=51540 29000 0 180 $X=50855 $Y=27485
X2595 94 32 37 333 31 444 447 NOR2_X1 $T=52110 26200 0 180 $X=51425 $Y=24685
X2596 62 32 142 334 31 444 448 NOR2_X1 $T=52110 26200 1 180 $X=51425 $Y=26085
X2597 332 32 335 337 31 443 446 NOR2_X1 $T=52110 23400 1 0 $X=51995 $Y=21885
X2598 61 32 95 63 31 240 448 NOR2_X1 $T=52110 29000 1 0 $X=51995 $Y=27485
X2599 336 32 18 261 31 445 446 NOR2_X1 $T=53440 20600 0 0 $X=53325 $Y=20485
X2600 262 32 337 392 31 443 447 NOR2_X1 $T=54580 23400 0 0 $X=54465 $Y=23285
X2601 20 32 96 413 31 445 241 NOR2_X1 $T=54770 20600 1 0 $X=54655 $Y=19085
X2602 301 32 413 412 31 445 446 NOR2_X1 $T=55910 20600 1 180 $X=55225 $Y=20485
X2603 97 32 98 265 31 445 241 NOR2_X1 $T=56860 20600 1 0 $X=56745 $Y=19085
X2604 343 32 265 394 31 445 446 NOR2_X1 $T=58190 20600 1 180 $X=57505 $Y=20485
X2605 414 32 413 302 31 445 446 NOR2_X1 $T=58190 20600 0 0 $X=58075 $Y=20485
X2606 60 32 105 264 31 443 447 NOR2_X1 $T=59520 23400 0 0 $X=59405 $Y=23285
X2607 347 32 23 266 31 445 241 NOR2_X1 $T=61040 20600 0 180 $X=60355 $Y=19085
X2608 91 32 99 346 31 444 447 NOR2_X1 $T=61420 26200 0 180 $X=60735 $Y=24685
X2609 62 32 22 416 31 444 447 NOR2_X1 $T=62560 26200 0 180 $X=61875 $Y=24685
X2610 102 32 101 349 31 240 448 NOR2_X1 $T=64270 29000 0 180 $X=63585 $Y=27485
X2611 103 32 147 351 31 240 448 NOR2_X1 $T=64840 29000 0 180 $X=64155 $Y=27485
X2612 169 32 65 396 31 444 448 NOR2_X1 $T=65410 26200 0 0 $X=65295 $Y=26085
X2613 68 32 274 352 31 445 446 NOR2_X1 $T=66740 20600 1 180 $X=66055 $Y=20485
X2614 60 32 65 277 31 444 448 NOR2_X1 $T=68450 26200 1 180 $X=67765 $Y=26085
X2615 91 32 105 427 31 444 447 NOR2_X1 $T=71490 26200 0 180 $X=70805 $Y=24685
X2616 62 32 99 375 31 240 448 NOR2_X1 $T=71680 29000 0 180 $X=70995 $Y=27485
X2617 92 32 22 171 31 240 448 NOR2_X1 $T=71680 29000 1 0 $X=71565 $Y=27485
X2618 279 32 355 106 31 445 241 NOR2_X1 $T=72060 20600 1 0 $X=71945 $Y=19085
X2619 102 32 150 398 31 443 446 NOR2_X1 $T=73770 23400 1 0 $X=73655 $Y=21885
X2620 428 32 106 357 31 445 446 NOR2_X1 $T=74720 20600 1 180 $X=74035 $Y=20485
X2621 103 32 54 358 31 443 446 NOR2_X1 $T=74340 23400 1 0 $X=74225 $Y=21885
X2622 26 32 13 108 31 240 448 NOR2_X1 $T=74910 29000 0 180 $X=74225 $Y=27485
X2623 50 32 150 304 31 444 448 NOR2_X1 $T=74530 26200 0 0 $X=74415 $Y=26085
X2624 94 32 85 135 31 240 448 NOR2_X1 $T=75480 29000 0 180 $X=74795 $Y=27485
X2625 169 32 55 376 31 443 447 NOR2_X1 $T=76620 23400 0 0 $X=76505 $Y=23285
X2626 417 32 282 112 31 445 241 NOR2_X1 $T=79280 20600 0 180 $X=78595 $Y=19085
X2627 60 32 145 429 31 444 448 NOR2_X1 $T=81180 26200 0 0 $X=81065 $Y=26085
X2628 92 32 105 185 31 240 448 NOR2_X1 $T=81180 29000 1 0 $X=81065 $Y=27485
X2629 91 32 101 402 31 443 447 NOR2_X1 $T=83460 23400 0 0 $X=83345 $Y=23285
X2630 62 32 147 403 31 444 447 NOR2_X1 $T=83460 26200 1 0 $X=83345 $Y=24685
X2631 94 32 22 173 31 240 448 NOR2_X1 $T=84790 29000 0 180 $X=84105 $Y=27485
X2632 31 412 371 263 32 443 446 XNOR2_X1 $T=54770 23400 1 0 $X=54655 $Y=21885
X2633 32 344 342 209 31 444 448 XOR2_X1 $T=54960 26200 0 0 $X=54845 $Y=26085
X2634 32 340 167 392 31 443 447 XOR2_X1 $T=55150 23400 0 0 $X=55035 $Y=23285
X2635 32 373 64 394 31 443 447 XOR2_X1 $T=56290 23400 0 0 $X=56175 $Y=23285
X2636 32 19 424 372 31 444 447 XOR2_X1 $T=56670 26200 1 0 $X=56555 $Y=24685
X2637 32 270 170 406 31 445 446 XOR2_X1 $T=70540 20600 1 180 $X=69285 $Y=20485
X2638 332 31 335 411 32 443 446 NAND2_X1 $T=51540 23400 1 0 $X=51425 $Y=21885
X2639 336 31 18 260 32 443 446 NAND2_X1 $T=53440 23400 1 0 $X=53325 $Y=21885
X2640 97 31 98 414 32 445 241 NAND2_X1 $T=58000 20600 0 180 $X=57315 $Y=19085
X2641 347 31 23 267 32 445 241 NAND2_X1 $T=61610 20600 0 180 $X=60925 $Y=19085
X2642 68 31 274 269 32 445 446 NAND2_X1 $T=68070 20600 0 0 $X=67955 $Y=20485
X2643 110 31 71 428 32 445 241 NAND2_X1 $T=74910 20600 1 0 $X=74795 $Y=19085
X2644 417 31 282 111 32 445 241 NAND2_X1 $T=78710 20600 0 180 $X=78025 $Y=19085
X2645 113 31 30 27 32 445 241 NAND2_X1 $T=83270 20600 0 180 $X=82585 $Y=19085
X2646 411 260 180 339 31 32 444 448 AOI21_X1 $T=53440 26200 0 0 $X=53325 $Y=26085
X2647 260 19 340 261 31 32 443 447 AOI21_X1 $T=53820 23400 0 0 $X=53705 $Y=23285
X2648 415 267 373 266 31 32 445 446 AOI21_X1 $T=60090 20600 0 0 $X=59975 $Y=20485
X2649 267 269 268 374 31 32 445 446 AOI21_X1 $T=60850 20600 0 0 $X=60735 $Y=20485
X2650 347 23 181 266 31 32 445 241 AOI21_X1 $T=62750 20600 0 180 $X=61875 $Y=19085
X2651 269 270 100 352 31 32 445 446 AOI21_X1 $T=64080 20600 1 180 $X=63205 $Y=20485
X2652 111 27 356 123 31 32 445 241 AOI21_X1 $T=78140 20600 0 180 $X=77265 $Y=19085
X2653 417 282 184 112 31 32 445 241 AOI21_X1 $T=80040 20600 0 180 $X=79165 $Y=19085
X2661 338 31 341 165 32 339 240 448 NAND3_X1 $T=54010 29000 1 0 $X=53895 $Y=27485
X2662 305 1 418 306 32 31 33 445 446 FA_X1 $T=1000 20600 0 0 $X=885 $Y=20485
X2663 430 305 72 407 32 31 73 443 446 FA_X1 $T=1000 23400 1 0 $X=885 $Y=21885
X2664 377 430 152 365 32 31 419 443 447 FA_X1 $T=1000 23400 0 0 $X=885 $Y=23285
X2665 126 419 198 309 32 31 378 444 448 FA_X1 $T=1000 26200 0 0 $X=885 $Y=26085
X2666 174 3 288 285 32 31 242 443 446 FA_X1 $T=4040 23400 1 0 $X=3925 $Y=21885
X2667 153 242 137 378 32 31 214 240 448 FA_X1 $T=7270 29000 0 180 $X=4115 $Y=27485
X2668 365 286 420 84 32 31 379 444 447 FA_X1 $T=9930 26200 0 180 $X=6775 $Y=24685
X2669 285 5 379 308 32 31 76 445 241 FA_X1 $T=7460 20600 1 0 $X=7345 $Y=19085
X2670 244 243 307 310 32 31 308 443 446 FA_X1 $T=7650 23400 1 0 $X=7535 $Y=21885
X2671 34 244 380 6 32 31 309 444 448 FA_X1 $T=8410 26200 0 0 $X=8295 $Y=26085
X2672 154 366 431 312 32 31 381 444 447 FA_X1 $T=9930 26200 1 0 $X=9815 $Y=24685
X2673 380 7 78 141 32 31 39 445 241 FA_X1 $T=10500 20600 1 0 $X=10385 $Y=19085
X2674 175 381 377 187 32 31 382 444 448 FA_X1 $T=11450 26200 0 0 $X=11335 $Y=26085
X2675 155 382 199 311 32 31 40 240 448 FA_X1 $T=11830 29000 1 0 $X=11715 $Y=27485
X2676 431 367 421 404 32 31 287 445 446 FA_X1 $T=12590 20600 0 0 $X=12475 $Y=20485
X2677 311 245 287 383 32 31 288 444 447 FA_X1 $T=12970 26200 1 0 $X=12855 $Y=24685
X2678 366 314 384 200 32 31 245 444 448 FA_X1 $T=14490 26200 0 0 $X=14375 $Y=26085
X2679 312 246 313 289 32 31 383 443 446 FA_X1 $T=14870 23400 1 0 $X=14755 $Y=21885
X2680 41 188 81 201 32 31 156 445 241 FA_X1 $T=16010 20600 1 0 $X=15895 $Y=19085
X2681 118 114 247 42 32 31 315 445 446 FA_X1 $T=18670 20600 0 0 $X=18555 $Y=20485
X2682 247 385 290 316 32 31 45 444 447 FA_X1 $T=21140 26200 1 0 $X=21025 $Y=24685
X2683 43 138 251 189 32 31 158 443 447 FA_X1 $T=21710 23400 0 0 $X=21595 $Y=23285
X2684 44 422 318 386 32 31 317 445 446 FA_X1 $T=23420 20600 0 0 $X=23305 $Y=20485
X2685 386 9 159 408 32 31 129 444 448 FA_X1 $T=25700 26200 0 0 $X=25585 $Y=26085
X2686 318 202 47 315 32 31 387 445 446 FA_X1 $T=26460 20600 0 0 $X=26345 $Y=20485
X2687 251 250 317 203 32 31 128 443 446 FA_X1 $T=30450 23400 0 180 $X=27295 $Y=21885
X2688 249 248 190 319 32 31 252 240 448 FA_X1 $T=27790 29000 1 0 $X=27675 $Y=27485
X2689 408 249 320 323 32 31 11 444 447 FA_X1 $T=28930 26200 1 0 $X=28815 $Y=24685
X2690 422 48 191 144 32 31 388 445 446 FA_X1 $T=29500 20600 0 0 $X=29385 $Y=20485
X2691 250 387 388 204 32 31 86 443 446 FA_X1 $T=30450 23400 1 0 $X=30335 $Y=21885
X2692 130 252 391 389 32 31 160 240 448 FA_X1 $T=30830 29000 1 0 $X=30715 $Y=27485
X2693 320 253 433 409 32 31 391 443 447 FA_X1 $T=33110 23400 0 0 $X=32995 $Y=23285
X2694 323 432 434 321 32 31 389 444 448 FA_X1 $T=36720 26200 1 180 $X=33565 $Y=26085
X2695 293 368 322 205 32 31 291 445 241 FA_X1 $T=38430 20600 0 180 $X=35275 $Y=19085
X2696 410 390 255 292 32 31 324 443 446 FA_X1 $T=35390 23400 1 0 $X=35275 $Y=21885
X2697 176 254 293 410 32 31 325 444 447 FA_X1 $T=35390 26200 1 0 $X=35275 $Y=24685
X2698 177 435 139 325 32 31 294 444 448 FA_X1 $T=36720 26200 0 0 $X=36605 $Y=26085
X2699 51 206 423 215 32 31 405 445 446 FA_X1 $T=38430 20600 0 0 $X=38315 $Y=20485
X2700 435 296 291 324 32 31 131 443 446 FA_X1 $T=41470 23400 0 180 $X=38315 $Y=21885
X2701 254 295 326 369 32 31 296 444 447 FA_X1 $T=38430 26200 1 0 $X=38315 $Y=24685
X2702 132 192 162 297 32 31 423 445 446 FA_X1 $T=41470 20600 0 0 $X=41355 $Y=20485
X2703 133 405 207 294 32 31 256 443 446 FA_X1 $T=41470 23400 1 0 $X=41355 $Y=21885
X2704 178 256 329 193 32 31 330 443 446 FA_X1 $T=44510 23400 1 0 $X=44395 $Y=21885
X2705 163 14 327 331 32 31 298 444 447 FA_X1 $T=45080 26200 1 0 $X=44965 $Y=24685
X2706 297 257 328 370 32 31 164 445 241 FA_X1 $T=45270 20600 1 0 $X=45155 $Y=19085
X2707 58 15 298 208 32 31 329 444 448 FA_X1 $T=45460 26200 0 0 $X=45345 $Y=26085
X2708 179 258 300 334 32 31 331 444 448 FA_X1 $T=48500 26200 0 0 $X=48385 $Y=26085
X2709 59 259 299 333 32 31 327 443 447 FA_X1 $T=48690 23400 0 0 $X=48575 $Y=23285
X2710 425 264 346 416 32 31 272 444 447 FA_X1 $T=57810 26200 1 0 $X=57695 $Y=24685
X2711 119 194 425 395 32 31 345 444 448 FA_X1 $T=61420 26200 1 180 $X=58265 $Y=26085
X2712 120 271 345 210 32 31 348 443 446 FA_X1 $T=64270 23400 0 180 $X=61115 $Y=21885
X2713 395 349 351 396 32 31 350 444 448 FA_X1 $T=61420 26200 0 0 $X=61305 $Y=26085
X2714 271 272 350 148 32 31 275 443 447 FA_X1 $T=63890 23400 0 0 $X=63775 $Y=23285
X2715 276 275 354 70 32 31 426 443 447 FA_X1 $T=66930 23400 0 0 $X=66815 $Y=23285
X2716 273 278 276 348 32 31 274 443 446 FA_X1 $T=70730 23400 0 180 $X=67575 $Y=21885
X2717 69 24 104 195 32 31 397 240 448 FA_X1 $T=68070 29000 1 0 $X=67955 $Y=27485
X2718 182 277 427 375 32 31 353 444 448 FA_X1 $T=68450 26200 0 0 $X=68335 $Y=26085
X2719 278 426 397 149 32 31 355 443 446 FA_X1 $T=70730 23400 1 0 $X=70615 $Y=21885
X2720 354 25 211 353 32 31 399 444 448 FA_X1 $T=71490 26200 0 0 $X=71375 $Y=26085
X2721 280 140 172 399 32 31 71 443 447 FA_X1 $T=73580 23400 0 0 $X=73465 $Y=23285
X2722 400 398 358 376 32 31 359 443 446 FA_X1 $T=78900 23400 0 180 $X=75745 $Y=21885
X2723 183 363 400 304 32 31 284 444 447 FA_X1 $T=77380 26200 1 0 $X=77265 $Y=24685
X2724 361 28 212 362 32 31 282 444 448 FA_X1 $T=78140 26200 0 0 $X=78025 $Y=26085
X2725 436 283 213 401 32 31 30 443 447 FA_X1 $T=80420 23400 0 0 $X=80305 $Y=23285
X2726 362 284 197 151 32 31 283 444 447 FA_X1 $T=80420 26200 1 0 $X=80305 $Y=24685
X2727 401 116 364 359 32 31 136 445 446 FA_X1 $T=81750 20600 0 0 $X=81635 $Y=20485
X2728 363 429 402 403 32 31 364 444 448 FA_X1 $T=81750 26200 0 0 $X=81635 $Y=26085
X2729 373 343 31 263 98 97 32 445 446 OAI22_X1 $T=55910 20600 0 0 $X=55795 $Y=20485
X2730 270 32 352 374 31 303 445 446 NOR3_X1 $T=63320 20600 1 180 $X=62445 $Y=20485
X2735 371 32 424 342 168 196 31 444 448 NOR4_X1 $T=57430 26200 0 0 $X=57315 $Y=26085
X2736 107 32 356 357 109 270 31 445 241 NOR4_X1 $T=73960 20600 1 0 $X=73845 $Y=19085
X2738 72 88 31 32 444 447 INV_X2 $T=5750 26200 1 0 $X=5635 $Y=24685
X2739 1 117 31 32 444 447 INV_X2 $T=6320 26200 1 0 $X=6205 $Y=24685
X2740 157 22 31 32 443 447 INV_X2 $T=20380 23400 0 0 $X=20265 $Y=23285
X2741 84 127 31 32 240 448 INV_X2 $T=20570 29000 1 0 $X=20455 $Y=27485
X2742 143 66 31 32 240 448 INV_X2 $T=21140 29000 1 0 $X=21025 $Y=27485
X2743 90 102 31 32 240 448 INV_X2 $T=35390 29000 1 0 $X=35275 $Y=27485
X2744 413 265 266 31 32 374 445 241 OR3_X1 $T=59520 20600 1 0 $X=59405 $Y=19085
.ENDS
***************************************
.SUBCKT ICV_18
** N=4 EP=0 IP=8 FDC=0
.ENDS
***************************************
.SUBCKT ICV_19 1 2 3 4 5 6 7 8 9 10 11 12 13 14 15 16 17 18 19 20
+ 21 22 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40
+ 41 42 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60
+ 61 62 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80
+ 81 82 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100
+ 101 102 103 104 105 106 107 108 109 110 111 112 113 114 115 116 117 118 119 120
+ 121 122 123 124 125 126 127 128 129 130 131 132 133 134 135 136 137 138 139 140
+ 141 142 143 144 145 146 147 148 149 150 151 152 153 154 155 156 157 158 159 160
+ 161 162 163 164 165 166 167 168 169 170 171 172 173 174 175 176 177 178 179 180
+ 181 182 183 184 185 186 187 188 189 190 191 192 193 194 195 196 197 198 199 200
+ 201 202 203 204 205 206 207 208 209 210 211 212 213 214 215 216 228 229
** N=463 EP=218 IP=5182 FDC=3078
X2429 349 284 23 24 91 458 463 AND2_X1 $T=83460 12200 1 0 $X=83345 $Y=10685
X2464 365 23 24 342 457 461 INV_X1 $T=78330 17800 0 180 $X=77835 $Y=16285
X2465 90 23 24 353 460 229 INV_X1 $T=84220 9400 0 180 $X=83725 $Y=7885
X2505 191 386 258 23 24 188 457 228 HA_X1 $T=54580 17800 0 0 $X=54465 $Y=17685
X2506 124 192 260 23 24 386 457 228 HA_X1 $T=58380 17800 1 180 $X=56365 $Y=17685
X2507 127 172 272 23 24 82 457 228 HA_X1 $T=69020 17800 0 0 $X=68905 $Y=17685
X2508 347 88 282 23 24 281 460 229 HA_X1 $T=82130 9400 0 180 $X=80115 $Y=7885
X2509 284 138 399 23 24 285 459 461 HA_X1 $T=84790 15000 1 180 $X=82775 $Y=14885
X2510 178 443 285 23 24 190 457 228 HA_X1 $T=82890 17800 0 0 $X=82775 $Y=17685
X2669 25 24 65 56 23 460 229 NOR2_X1 $T=5560 9400 1 0 $X=5445 $Y=7885
X2670 30 24 48 103 23 458 462 NOR2_X1 $T=5750 12200 0 0 $X=5635 $Y=12085
X2671 5 24 35 57 23 460 463 NOR2_X1 $T=8600 9400 0 0 $X=8485 $Y=9285
X2672 5 24 58 233 23 459 462 NOR2_X1 $T=9550 15000 0 180 $X=8865 $Y=13485
X2673 151 24 94 419 23 459 461 NOR2_X1 $T=9550 15000 1 180 $X=8865 $Y=14885
X2674 45 24 68 420 23 457 461 NOR2_X1 $T=9740 17800 0 180 $X=9055 $Y=16285
X2675 27 24 37 371 23 459 461 NOR2_X1 $T=11070 15000 1 180 $X=10385 $Y=14885
X2676 25 24 58 158 23 457 228 NOR2_X1 $T=10500 17800 0 0 $X=10385 $Y=17685
X2677 141 24 26 401 23 458 462 NOR2_X1 $T=11260 12200 1 180 $X=10575 $Y=12085
X2678 28 24 12 299 23 459 462 NOR2_X1 $T=11640 15000 1 0 $X=11525 $Y=13485
X2679 74 24 29 234 23 459 461 NOR2_X1 $T=12020 15000 0 0 $X=11905 $Y=14885
X2680 61 24 29 235 23 458 462 NOR2_X1 $T=13540 12200 1 180 $X=12855 $Y=12085
X2681 5 24 12 160 23 457 228 NOR2_X1 $T=13540 17800 1 180 $X=12855 $Y=17685
X2682 28 24 26 161 23 457 228 NOR2_X1 $T=14110 17800 1 180 $X=13425 $Y=17685
X2683 61 24 142 300 23 457 461 NOR2_X1 $T=14870 17800 0 180 $X=14185 $Y=16285
X2684 25 24 48 162 23 460 229 NOR2_X1 $T=15060 9400 1 0 $X=14945 $Y=7885
X2685 5 24 65 106 23 460 463 NOR2_X1 $T=16770 9400 1 180 $X=16085 $Y=9285
X2686 28 24 35 95 23 460 229 NOR2_X1 $T=17150 9400 0 180 $X=16465 $Y=7885
X2687 30 24 34 447 23 459 462 NOR2_X1 $T=18100 15000 0 180 $X=17415 $Y=13485
X2688 5 24 48 163 23 460 463 NOR2_X1 $T=18860 9400 0 0 $X=18745 $Y=9285
X2689 30 24 78 423 23 459 461 NOR2_X1 $T=19050 15000 0 0 $X=18935 $Y=14885
X2690 28 24 65 64 23 460 229 NOR2_X1 $T=19430 9400 1 0 $X=19315 $Y=7885
X2691 25 24 34 402 23 457 461 NOR2_X1 $T=19810 17800 1 0 $X=19695 $Y=16285
X2692 32 24 142 355 23 458 462 NOR2_X1 $T=20190 12200 0 0 $X=20075 $Y=12085
X2693 141 24 35 96 23 460 463 NOR2_X1 $T=20760 9400 0 0 $X=20645 $Y=9285
X2694 32 24 29 240 23 458 463 NOR2_X1 $T=22850 12200 1 0 $X=22735 $Y=10685
X2695 30 24 42 241 23 459 462 NOR2_X1 $T=23800 15000 1 0 $X=23685 $Y=13485
X2696 5 24 34 426 23 458 462 NOR2_X1 $T=26080 12200 1 180 $X=25395 $Y=12085
X2697 25 24 78 427 23 459 461 NOR2_X1 $T=26270 15000 1 180 $X=25585 $Y=14885
X2698 141 24 48 448 23 457 461 NOR2_X1 $T=26840 17800 1 0 $X=26725 $Y=16285
X2699 36 24 142 425 23 460 229 NOR2_X1 $T=27790 9400 0 180 $X=27105 $Y=7885
X2700 36 24 29 303 23 458 463 NOR2_X1 $T=27410 12200 1 0 $X=27295 $Y=10685
X2701 45 24 65 377 23 457 228 NOR2_X1 $T=27410 17800 0 0 $X=27295 $Y=17685
X2702 151 24 35 428 23 459 461 NOR2_X1 $T=28170 15000 0 0 $X=28055 $Y=14885
X2703 61 24 68 165 23 460 229 NOR2_X1 $T=30070 9400 1 0 $X=29955 $Y=7885
X2704 144 24 142 429 23 460 463 NOR2_X1 $T=30070 9400 0 0 $X=29955 $Y=9285
X2705 27 24 58 245 23 460 463 NOR2_X1 $T=30640 9400 0 0 $X=30525 $Y=9285
X2706 36 24 37 69 23 460 463 NOR2_X1 $T=31210 9400 0 0 $X=31095 $Y=9285
X2707 61 24 26 244 23 458 463 NOR2_X1 $T=31780 12200 1 0 $X=31665 $Y=10685
X2708 32 24 68 246 23 459 462 NOR2_X1 $T=31970 15000 1 0 $X=31855 $Y=13485
X2709 74 24 12 430 23 458 463 NOR2_X1 $T=32350 12200 1 0 $X=32235 $Y=10685
X2710 36 24 94 306 23 457 461 NOR2_X1 $T=34060 17800 0 180 $X=33375 $Y=16285
X2711 144 24 37 449 23 459 462 NOR2_X1 $T=34060 15000 1 0 $X=33945 $Y=13485
X2712 144 24 29 243 23 457 228 NOR2_X1 $T=34630 17800 1 180 $X=33945 $Y=17685
X2713 145 24 38 248 23 458 462 NOR2_X1 $T=34820 12200 0 0 $X=34705 $Y=12085
X2714 61 24 147 308 23 457 461 NOR2_X1 $T=36150 17800 1 0 $X=36035 $Y=16285
X2715 72 24 40 73 23 460 463 NOR2_X1 $T=36340 9400 0 0 $X=36225 $Y=9285
X2716 32 24 41 405 23 459 462 NOR2_X1 $T=36340 15000 1 0 $X=36225 $Y=13485
X2717 149 24 42 357 23 458 462 NOR2_X1 $T=36530 12200 0 0 $X=36415 $Y=12085
X2718 39 24 34 168 23 457 228 NOR2_X1 $T=36530 17800 0 0 $X=36415 $Y=17685
X2719 74 24 148 247 23 457 461 NOR2_X1 $T=36720 17800 1 0 $X=36605 $Y=16285
X2720 145 24 40 249 23 460 463 NOR2_X1 $T=38430 9400 1 180 $X=37745 $Y=9285
X2721 39 24 78 358 23 458 462 NOR2_X1 $T=38050 12200 0 0 $X=37935 $Y=12085
X2722 45 24 15 450 23 457 461 NOR2_X1 $T=38620 17800 1 0 $X=38505 $Y=16285
X2723 27 24 87 406 23 459 461 NOR2_X1 $T=39570 15000 0 0 $X=39455 $Y=14885
X2724 149 24 38 309 23 458 463 NOR2_X1 $T=39760 12200 1 0 $X=39645 $Y=10685
X2725 39 24 42 310 23 460 463 NOR2_X1 $T=40140 9400 0 0 $X=40025 $Y=9285
X2726 151 24 52 451 23 457 461 NOR2_X1 $T=41090 17800 0 180 $X=40405 $Y=16285
X2727 46 24 34 253 23 459 461 NOR2_X1 $T=41660 15000 0 0 $X=41545 $Y=14885
X2728 46 24 78 251 23 460 463 NOR2_X1 $T=42610 9400 0 0 $X=42495 $Y=9285
X2729 10 24 34 290 23 458 463 NOR2_X1 $T=44130 12200 0 180 $X=43445 $Y=10685
X2730 10 24 48 381 23 459 462 NOR2_X1 $T=44320 15000 1 0 $X=44205 $Y=13485
X2731 11 24 48 359 23 460 463 NOR2_X1 $T=45650 9400 1 180 $X=44965 $Y=9285
X2732 11 24 65 382 23 459 461 NOR2_X1 $T=46410 15000 1 180 $X=45725 $Y=14885
X2733 53 24 35 316 23 460 463 NOR2_X1 $T=46220 9400 0 0 $X=46105 $Y=9285
X2734 76 24 58 432 23 458 463 NOR2_X1 $T=48690 12200 0 180 $X=48005 $Y=10685
X2735 77 24 12 409 23 458 463 NOR2_X1 $T=49260 12200 0 180 $X=48575 $Y=10685
X2736 145 24 44 255 23 460 463 NOR2_X1 $T=52490 9400 0 0 $X=52375 $Y=9285
X2737 149 24 40 320 23 458 463 NOR2_X1 $T=54010 12200 1 0 $X=53895 $Y=10685
X2738 39 24 38 361 23 460 463 NOR2_X1 $T=55530 9400 1 180 $X=54845 $Y=9285
X2739 46 24 42 256 23 460 463 NOR2_X1 $T=55530 9400 0 0 $X=55415 $Y=9285
X2740 11 24 34 387 23 458 462 NOR2_X1 $T=58000 12200 1 180 $X=57315 $Y=12085
X2741 10 24 78 322 23 458 463 NOR2_X1 $T=58190 12200 0 180 $X=57505 $Y=10685
X2742 36 24 87 263 23 458 462 NOR2_X1 $T=60090 12200 0 0 $X=59975 $Y=12085
X2743 144 24 148 329 23 458 463 NOR2_X1 $T=60280 12200 1 0 $X=60165 $Y=10685
X2744 46 24 38 388 23 460 463 NOR2_X1 $T=60660 9400 0 0 $X=60545 $Y=9285
X2745 72 24 147 412 23 458 462 NOR2_X1 $T=62370 12200 0 0 $X=62255 $Y=12085
X2746 10 24 42 325 23 460 463 NOR2_X1 $T=63320 9400 1 180 $X=62635 $Y=9285
X2747 11 24 78 328 23 460 229 NOR2_X1 $T=63510 9400 0 180 $X=62825 $Y=7885
X2748 61 24 15 436 23 458 462 NOR2_X1 $T=64270 12200 0 0 $X=64155 $Y=12085
X2749 145 24 41 267 23 460 229 NOR2_X1 $T=64650 9400 1 0 $X=64535 $Y=7885
X2750 32 24 52 390 23 459 461 NOR2_X1 $T=65220 15000 0 0 $X=65105 $Y=14885
X2751 149 24 44 332 23 458 463 NOR2_X1 $T=67500 12200 0 180 $X=66815 $Y=10685
X2752 36 24 52 293 23 459 461 NOR2_X1 $T=67500 15000 1 180 $X=66815 $Y=14885
X2753 39 24 40 333 23 460 463 NOR2_X1 $T=67880 9400 1 180 $X=67195 $Y=9285
X2754 53 24 34 270 23 459 462 NOR2_X1 $T=68070 15000 0 180 $X=67385 $Y=13485
X2755 144 24 87 334 23 457 228 NOR2_X1 $T=68450 17800 0 0 $X=68335 $Y=17685
X2756 10 24 15 81 23 458 463 NOR2_X1 $T=68640 12200 1 0 $X=68525 $Y=10685
X2757 11 24 52 171 23 460 229 NOR2_X1 $T=69400 9400 0 180 $X=68715 $Y=7885
X2758 77 24 65 363 23 459 462 NOR2_X1 $T=69590 15000 0 180 $X=68905 $Y=13485
X2759 76 24 48 438 23 458 463 NOR2_X1 $T=69780 12200 0 180 $X=69095 $Y=10685
X2760 72 24 148 413 23 459 461 NOR2_X1 $T=69210 15000 0 0 $X=69095 $Y=14885
X2761 46 24 15 271 23 458 463 NOR2_X1 $T=69780 12200 1 0 $X=69665 $Y=10685
X2762 149 24 15 440 23 458 463 NOR2_X1 $T=71490 12200 0 180 $X=70805 $Y=10685
X2763 10 24 52 364 23 460 463 NOR2_X1 $T=71110 9400 0 0 $X=70995 $Y=9285
X2764 11 24 87 391 23 460 463 NOR2_X1 $T=71680 9400 0 0 $X=71565 $Y=9285
X2765 173 24 55 337 23 457 228 NOR2_X1 $T=72060 17800 0 0 $X=71945 $Y=17685
X2766 39 24 52 414 23 458 463 NOR2_X1 $T=73200 12200 0 180 $X=72515 $Y=10685
X2767 39 24 15 86 23 460 463 NOR2_X1 $T=73960 9400 0 0 $X=73845 $Y=9285
X2768 46 24 52 277 23 460 463 NOR2_X1 $T=74530 9400 0 0 $X=74415 $Y=9285
X2769 85 24 276 441 23 457 461 NOR2_X1 $T=74720 17800 1 0 $X=74605 $Y=16285
X2770 176 24 175 276 23 457 228 NOR2_X1 $T=74720 17800 0 0 $X=74605 $Y=17685
X2771 46 24 87 295 23 457 461 NOR2_X1 $T=75290 17800 1 0 $X=75175 $Y=16285
X2772 10 24 87 345 23 458 462 NOR2_X1 $T=76050 12200 1 180 $X=75365 $Y=12085
X2773 10 24 148 343 23 458 462 NOR2_X1 $T=76050 12200 0 0 $X=75935 $Y=12085
X2774 11 24 147 341 23 457 461 NOR2_X1 $T=76620 17800 1 0 $X=76505 $Y=16285
X2775 11 24 148 392 23 458 462 NOR2_X1 $T=78140 12200 1 180 $X=77455 $Y=12085
X2776 53 24 41 280 23 459 462 NOR2_X1 $T=78900 15000 1 0 $X=78785 $Y=13485
X2777 76 24 44 346 23 457 461 NOR2_X1 $T=80230 17800 1 0 $X=80115 $Y=16285
X2778 77 24 40 394 23 459 461 NOR2_X1 $T=81750 15000 1 180 $X=81065 $Y=14885
X2779 347 24 283 89 23 460 229 NOR2_X1 $T=82130 9400 1 0 $X=82015 $Y=7885
X2780 178 24 177 278 23 457 228 NOR2_X1 $T=82890 17800 1 180 $X=82205 $Y=17685
X2781 353 24 89 398 23 460 229 NOR2_X1 $T=83270 9400 0 180 $X=82585 $Y=7885
X2782 284 24 349 92 23 458 463 NOR2_X1 $T=82890 12200 1 0 $X=82775 $Y=10685
X2783 91 24 92 416 23 458 463 NOR2_X1 $T=84790 12200 0 180 $X=84105 $Y=10685
X2784 23 337 335 273 24 457 228 XNOR2_X1 $T=72060 17800 1 180 $X=70805 $Y=17685
X2785 23 416 351 444 24 459 462 XNOR2_X1 $T=84790 15000 0 180 $X=83535 $Y=13485
X2786 24 125 326 199 23 457 228 XOR2_X1 $T=63700 17800 1 180 $X=62445 $Y=17685
X2787 24 294 336 441 23 457 461 XOR2_X1 $T=74720 17800 0 180 $X=73465 $Y=16285
X2788 24 365 415 131 23 457 461 XOR2_X1 $T=79090 17800 1 0 $X=78975 $Y=16285
X2789 24 132 352 398 23 460 463 XOR2_X1 $T=82130 9400 1 180 $X=80875 $Y=9285
X2790 24 19 350 202 23 457 461 XOR2_X1 $T=81940 17800 1 0 $X=81825 $Y=16285
X2791 347 23 283 90 24 460 229 NAND2_X1 $T=84790 9400 0 180 $X=84105 $Y=7885
X2792 342 17 294 16 23 24 457 461 AOI21_X1 $T=77950 17800 0 180 $X=77075 $Y=16285
X2793 189 19 365 278 23 24 457 228 AOI21_X1 $T=80230 17800 1 180 $X=79355 $Y=17685
X2796 395 230 156 369 24 23 236 460 463 FA_X1 $T=1000 9400 0 0 $X=885 $Y=9285
X2797 21 1 417 354 24 23 366 458 462 FA_X1 $T=1000 12200 0 0 $X=885 $Y=12085
X2798 179 446 367 139 24 23 231 457 461 FA_X1 $T=1000 17800 1 0 $X=885 $Y=16285
X2799 417 2 296 400 24 23 368 458 463 FA_X1 $T=4040 12200 1 0 $X=3925 $Y=10685
X2800 418 420 419 371 24 23 297 459 461 FA_X1 $T=5940 15000 0 0 $X=5825 $Y=14885
X2801 445 233 299 401 24 23 370 458 462 FA_X1 $T=6320 12200 0 0 $X=6205 $Y=12085
X2802 446 193 421 368 24 23 298 458 463 FA_X1 $T=10120 12200 0 180 $X=6965 $Y=10685
X2803 230 3 194 205 24 23 59 460 229 FA_X1 $T=7840 9400 1 0 $X=7725 $Y=7885
X2804 400 235 355 140 24 23 105 458 463 FA_X1 $T=13160 12200 0 180 $X=10005 $Y=10685
X2805 232 234 300 182 24 23 372 457 461 FA_X1 $T=10690 17800 1 0 $X=10575 $Y=16285
X2806 296 4 60 33 24 23 373 460 229 FA_X1 $T=10880 9400 1 0 $X=10765 $Y=7885
X2807 159 236 396 298 24 23 62 459 462 FA_X1 $T=12210 15000 1 0 $X=12095 $Y=13485
X2808 215 374 63 447 24 23 375 459 461 FA_X1 $T=12590 15000 0 0 $X=12475 $Y=14885
X2809 396 206 422 238 24 23 107 458 462 FA_X1 $T=13540 12200 0 0 $X=13425 $Y=12085
X2810 374 195 423 402 24 23 301 457 228 FA_X1 $T=14110 17800 0 0 $X=13995 $Y=17685
X2811 238 424 302 287 24 23 286 459 462 FA_X1 $T=18100 15000 1 0 $X=17985 $Y=13485
X2812 31 239 286 7 24 23 110 457 228 FA_X1 $T=20190 17800 0 0 $X=20075 $Y=17685
X2813 239 134 397 376 24 23 111 457 461 FA_X1 $T=20380 17800 1 0 $X=20265 $Y=16285
X2814 108 240 425 70 24 23 66 460 463 FA_X1 $T=21330 9400 0 0 $X=21215 $Y=9285
X2815 287 242 209 208 24 23 376 458 463 FA_X1 $T=24370 12200 1 0 $X=24255 $Y=10685
X2816 97 304 288 143 24 23 67 460 463 FA_X1 $T=27030 9400 0 0 $X=26915 $Y=9285
X2817 378 303 429 71 24 23 242 458 463 FA_X1 $T=28740 12200 1 0 $X=28625 $Y=10685
X2818 304 8 289 404 24 23 114 459 462 FA_X1 $T=28930 15000 1 0 $X=28815 $Y=13485
X2819 9 307 305 403 24 23 113 457 461 FA_X1 $T=33490 17800 0 180 $X=30335 $Y=16285
X2820 404 245 430 244 24 23 305 458 462 FA_X1 $T=31780 12200 0 0 $X=31665 $Y=12085
X2821 183 356 167 146 24 23 407 460 463 FA_X1 $T=33300 9400 0 0 $X=33185 $Y=9285
X2822 289 246 306 449 24 23 307 459 461 FA_X1 $T=33490 15000 0 0 $X=33375 $Y=14885
X2823 116 247 308 405 24 23 250 459 461 FA_X1 $T=36530 15000 0 0 $X=36415 $Y=14885
X2824 356 248 357 358 24 23 408 458 463 FA_X1 $T=36720 12200 1 0 $X=36605 $Y=10685
X2825 184 196 312 407 24 23 379 458 462 FA_X1 $T=38620 12200 0 0 $X=38505 $Y=12085
X2826 47 135 314 452 24 23 254 457 461 FA_X1 $T=42040 17800 1 0 $X=41925 $Y=16285
X2827 185 254 291 152 24 23 317 457 228 FA_X1 $T=44130 17800 0 0 $X=44015 $Y=17685
X2828 453 456 315 383 24 23 431 459 462 FA_X1 $T=47930 15000 0 180 $X=44775 $Y=13485
X2829 75 453 379 317 24 23 433 459 461 FA_X1 $T=46410 15000 0 0 $X=46295 $Y=14885
X2830 186 433 313 99 24 23 120 457 228 FA_X1 $T=47170 17800 0 0 $X=47055 $Y=17685
X2831 291 198 360 197 24 23 383 460 463 FA_X1 $T=49450 9400 0 0 $X=49335 $Y=9285
X2832 187 13 454 431 24 23 121 457 461 FA_X1 $T=49830 17800 1 0 $X=49715 $Y=16285
X2833 315 212 434 385 24 23 384 458 462 FA_X1 $T=50400 12200 0 0 $X=50285 $Y=12085
X2834 360 137 319 292 24 23 434 458 463 FA_X1 $T=50970 12200 1 0 $X=50855 $Y=10685
X2835 292 255 320 361 24 23 49 460 229 FA_X1 $T=51920 9400 1 0 $X=51805 $Y=7885
X2836 258 257 213 323 24 23 122 457 461 FA_X1 $T=55910 17800 0 180 $X=52755 $Y=16285
X2837 454 384 321 203 24 23 257 459 462 FA_X1 $T=53250 15000 1 0 $X=53135 $Y=13485
X2838 319 256 322 387 24 23 123 458 463 FA_X1 $T=54580 12200 1 0 $X=54465 $Y=10685
X2839 50 261 435 410 24 23 79 460 463 FA_X1 $T=57620 9400 0 0 $X=57505 $Y=9285
X2840 261 388 325 328 24 23 327 460 229 FA_X1 $T=59900 9400 1 0 $X=59785 $Y=7885
X2841 259 265 436 390 24 23 330 459 462 FA_X1 $T=62370 15000 1 0 $X=62255 $Y=13485
X2842 435 267 332 333 24 23 331 460 463 FA_X1 $T=64270 9400 0 0 $X=64155 $Y=9285
X2843 324 268 330 154 24 23 269 457 461 FA_X1 $T=64460 17800 1 0 $X=64345 $Y=16285
X2844 455 270 438 363 24 23 266 458 462 FA_X1 $T=67880 12200 1 180 $X=64725 $Y=12085
X2845 362 269 437 155 24 23 272 457 228 FA_X1 $T=65410 17800 0 0 $X=65295 $Y=17685
X2846 265 293 334 413 24 23 128 457 461 FA_X1 $T=67500 17800 1 0 $X=67385 $Y=16285
X2847 100 271 364 391 24 23 101 460 229 FA_X1 $T=69400 9400 1 0 $X=69285 $Y=7885
X2848 274 275 440 414 24 23 279 458 462 FA_X1 $T=75480 12200 1 180 $X=72325 $Y=12085
X2849 348 279 201 214 24 23 282 460 463 FA_X1 $T=77950 9400 0 0 $X=77835 $Y=9285
X2850 339 280 346 394 24 23 393 459 461 FA_X1 $T=78140 15000 0 0 $X=78025 $Y=14885
X2851 399 20 393 344 24 23 283 458 462 FA_X1 $T=81750 12200 0 0 $X=81635 $Y=12085
X2852 294 85 23 273 175 176 24 457 228 OAI22_X1 $T=73770 17800 0 0 $X=73655 $Y=17685
X2853 132 353 23 444 283 347 24 460 463 OAI22_X1 $T=83840 9400 0 0 $X=83725 $Y=9285
X2854 19 24 278 18 23 200 457 228 NOR3_X1 $T=78140 17800 1 180 $X=77265 $Y=17685
X2859 22 231 395 366 24 23 102 354 372 297 370 369 459 462 ICV_9 $T=1000 15000 1 0 $X=885 $Y=13485
X2860 180 204 157 93 24 23 367 181 232 418 445 104 457 228 ICV_9 $T=1000 17800 0 0 $X=885 $Y=17685
X2861 421 237 133 373 24 23 422 237 375 216 378 424 458 463 ICV_9 $T=13160 12200 1 0 $X=13045 $Y=10685
X2862 302 6 301 207 24 23 397 109 241 427 426 164 459 461 ICV_9 $T=19620 15000 0 0 $X=19505 $Y=14885
X2863 112 448 377 428 24 23 403 288 243 166 210 115 457 228 ICV_9 $T=27980 17800 0 0 $X=27865 $Y=17685
X2864 169 249 309 310 24 23 170 98 251 290 359 119 460 229 ICV_9 $T=37860 9400 1 0 $X=37745 $Y=7885
X2865 43 450 451 406 24 23 311 118 252 136 211 313 457 228 ICV_9 $T=38050 17800 0 0 $X=37935 $Y=17685
X2866 117 250 311 150 24 23 252 452 253 381 382 380 459 462 ICV_9 $T=38240 15000 1 0 $X=38125 $Y=13485
X2867 312 318 380 408 24 23 456 314 316 432 409 318 458 462 ICV_9 $T=41660 12200 0 0 $X=41545 $Y=12085
X2868 385 259 51 455 24 23 262 321 262 324 411 389 459 462 ICV_9 $T=56290 15000 1 0 $X=56175 $Y=13485
X2869 323 14 80 153 24 23 264 260 264 362 389 126 457 461 ICV_9 $T=58380 17800 1 0 $X=58265 $Y=16285
X2870 410 263 329 412 24 23 268 411 266 327 331 437 458 463 ICV_9 $T=60850 12200 1 0 $X=60735 $Y=10685
X2871 129 274 339 340 24 23 442 340 295 343 341 344 459 462 ICV_9 $T=72820 15000 1 0 $X=72705 $Y=13485
X2872 275 277 345 392 24 23 130 443 281 348 442 349 458 463 ICV_9 $T=76810 12200 1 0 $X=76695 $Y=10685
X2875 336 24 335 83 326 439 23 457 461 NOR4_X1 $T=71490 17800 0 180 $X=70425 $Y=16285
X2876 352 24 351 350 415 338 23 459 462 NOR4_X1 $T=83650 15000 0 180 $X=82585 $Y=13485
X2877 54 23 84 439 338 174 24 459 462 NAND4_X1 $T=71870 15000 1 0 $X=71755 $Y=13485
X2878 63 78 23 24 457 461 INV_X2 $T=16200 17800 1 0 $X=16085 $Y=16285
X2879 33 34 23 24 458 462 INV_X2 $T=22660 12200 0 0 $X=22545 $Y=12085
X2880 70 144 23 24 457 461 INV_X2 $T=34060 17800 1 0 $X=33945 $Y=16285
X2881 71 72 23 24 459 462 INV_X2 $T=34630 15000 1 0 $X=34515 $Y=13485
X2882 140 36 23 24 457 228 INV_X2 $T=34630 17800 0 0 $X=34515 $Y=17685
X2883 55 276 16 23 24 18 457 228 OR3_X1 $T=76430 17800 0 0 $X=76315 $Y=17685
.ENDS
***************************************
.SUBCKT ICV_20 1 2 3 4 5 6 7 8 9 10 11 12 13 14 16 18 19 20 21 22
+ 23 24 25 26 27 28 29 30 31 32 33 34 35 36 37 38 39 40 41 42
+ 43 44 45 46 47 48 49 50 51 52 53 54 55 56 57 58 59 60 61 62
+ 63 64 65 66 67 68 69 70 71 72 73 74 75 76 77 78 79 80 81 82
+ 83 84 85 86 87 88 89 90 91 92 93 94 95 96 97 98 99 100 101 102
+ 103 104 105 106 107 108 109 110 111 112 113 114 115 122
** N=301 EP=114 IP=3599 FDC=2002
X1726 261 163 8 9 222 297 300 AND2_X1 $T=73580 1000 0 0 $X=73465 $Y=885
X1742 179 154 212 156 8 9 298 301 OAI21_X1 $T=60660 6600 1 0 $X=60545 $Y=5085
X1743 180 155 259 213 8 9 299 300 OAI21_X1 $T=62940 3800 1 0 $X=62825 $Y=2285
X1744 216 158 217 215 8 9 297 300 OAI21_X1 $T=66170 1000 0 0 $X=66055 $Y=885
X1745 216 158 240 218 8 9 299 300 OAI21_X1 $T=66170 3800 1 0 $X=66055 $Y=2285
X1746 267 165 266 173 8 9 297 300 OAI21_X1 $T=75860 1000 0 0 $X=75745 $Y=885
X1747 212 8 9 292 298 122 INV_X1 $T=61230 6600 0 0 $X=61115 $Y=6485
X1748 229 8 9 283 299 300 INV_X1 $T=80420 3800 1 0 $X=80305 $Y=2285
X1765 155 214 157 8 9 219 299 301 HA_X1 $T=63700 3800 0 0 $X=63585 $Y=3685
X1766 216 219 159 8 9 160 298 301 HA_X1 $T=65980 6600 1 0 $X=65865 $Y=5085
X1767 163 220 161 8 9 294 299 300 HA_X1 $T=70350 3800 0 180 $X=68335 $Y=2285
X1768 267 294 167 8 9 168 299 300 HA_X1 $T=76810 3800 1 0 $X=76695 $Y=2285
X1769 228 265 168 8 9 38 299 301 HA_X1 $T=79280 3800 1 180 $X=77265 $Y=3685
X1863 26 9 61 126 8 297 300 NOR2_X1 $T=9170 1000 1 180 $X=8485 $Y=885
X1864 16 9 76 232 8 299 301 NOR2_X1 $T=8790 3800 0 0 $X=8675 $Y=3685
X1865 10 9 25 270 8 299 301 NOR2_X1 $T=9930 3800 1 180 $X=9245 $Y=3685
X1866 68 9 59 246 8 299 301 NOR2_X1 $T=9930 3800 0 0 $X=9815 $Y=3685
X1867 28 9 24 125 8 299 301 NOR2_X1 $T=10500 3800 0 0 $X=10385 $Y=3685
X1868 14 9 60 185 8 299 300 NOR2_X1 $T=11260 3800 1 0 $X=11145 $Y=2285
X1869 68 9 24 285 8 298 122 NOR2_X1 $T=12780 6600 0 0 $X=12665 $Y=6485
X1870 10 9 59 286 8 299 301 NOR2_X1 $T=13540 3800 1 180 $X=12855 $Y=3685
X1871 16 9 61 129 8 299 300 NOR2_X1 $T=13730 3800 1 0 $X=13615 $Y=2285
X1872 26 9 25 271 8 299 301 NOR2_X1 $T=15440 3800 1 180 $X=14755 $Y=3685
X1873 13 9 60 189 8 299 300 NOR2_X1 $T=16770 3800 0 180 $X=16085 $Y=2285
X1874 14 9 76 233 8 299 301 NOR2_X1 $T=17340 3800 1 180 $X=16655 $Y=3685
X1875 14 9 61 132 8 299 301 NOR2_X1 $T=19430 3800 0 0 $X=19315 $Y=3685
X1876 13 9 76 191 8 299 301 NOR2_X1 $T=22850 3800 1 180 $X=22165 $Y=3685
X1877 12 9 60 274 8 297 300 NOR2_X1 $T=23040 1000 1 180 $X=22355 $Y=885
X1878 10 9 24 133 8 299 300 NOR2_X1 $T=24370 3800 1 0 $X=24255 $Y=2285
X1879 26 9 59 251 8 297 300 NOR2_X1 $T=26650 1000 1 180 $X=25965 $Y=885
X1880 16 9 25 192 8 299 300 NOR2_X1 $T=27790 3800 0 180 $X=27105 $Y=2285
X1881 26 9 24 135 8 299 300 NOR2_X1 $T=28550 3800 1 0 $X=28435 $Y=2285
X1882 28 9 67 137 8 298 301 NOR2_X1 $T=31590 6600 1 0 $X=31475 $Y=5085
X1883 14 9 25 195 8 297 300 NOR2_X1 $T=32350 1000 0 0 $X=32235 $Y=885
X1884 12 9 76 288 8 298 122 NOR2_X1 $T=32920 6600 1 180 $X=32235 $Y=6485
X1885 16 9 59 287 8 297 300 NOR2_X1 $T=32920 1000 0 0 $X=32805 $Y=885
X1886 68 9 35 289 8 298 301 NOR2_X1 $T=33490 6600 0 180 $X=32805 $Y=5085
X1887 10 9 3 275 8 298 301 NOR2_X1 $T=34060 6600 0 180 $X=33375 $Y=5085
X1888 29 9 37 138 8 298 122 NOR2_X1 $T=34440 6600 1 180 $X=33755 $Y=6485
X1889 12 9 30 196 8 297 300 NOR2_X1 $T=34630 1000 0 0 $X=34515 $Y=885
X1890 29 9 30 140 8 298 301 NOR2_X1 $T=35200 6600 1 0 $X=35085 $Y=5085
X1891 31 9 4 177 8 298 301 NOR2_X1 $T=35770 6600 1 0 $X=35655 $Y=5085
X1892 13 9 69 197 8 299 300 NOR2_X1 $T=36910 3800 1 0 $X=36795 $Y=2285
X1893 31 9 37 198 8 298 301 NOR2_X1 $T=37100 6600 1 0 $X=36985 $Y=5085
X1894 14 9 19 139 8 297 300 NOR2_X1 $T=38810 1000 1 180 $X=38125 $Y=885
X1895 33 9 4 199 8 298 301 NOR2_X1 $T=39000 6600 0 180 $X=38315 $Y=5085
X1896 26 9 18 200 8 299 300 NOR2_X1 $T=39950 3800 1 0 $X=39835 $Y=2285
X1897 16 9 34 202 8 299 300 NOR2_X1 $T=41850 3800 1 0 $X=41735 $Y=2285
X1898 14 9 34 145 8 299 300 NOR2_X1 $T=44510 3800 0 180 $X=43825 $Y=2285
X1899 12 9 69 205 8 299 300 NOR2_X1 $T=46600 3800 0 180 $X=45915 $Y=2285
X1900 13 9 19 255 8 297 300 NOR2_X1 $T=47170 1000 1 180 $X=46485 $Y=885
X1901 21 9 35 147 8 299 301 NOR2_X1 $T=47930 3800 0 0 $X=47815 $Y=3685
X1902 16 9 18 277 8 297 300 NOR2_X1 $T=48310 1000 0 0 $X=48195 $Y=885
X1903 36 9 24 278 8 299 301 NOR2_X1 $T=50210 3800 1 180 $X=49525 $Y=3685
X1904 20 9 3 207 8 298 301 NOR2_X1 $T=50590 6600 0 180 $X=49905 $Y=5085
X1905 29 9 69 234 8 299 301 NOR2_X1 $T=51540 3800 0 0 $X=51425 $Y=3685
X1906 31 9 30 235 8 299 301 NOR2_X1 $T=52110 3800 0 0 $X=51995 $Y=3685
X1907 33 9 37 236 8 299 301 NOR2_X1 $T=52680 3800 0 0 $X=52565 $Y=3685
X1908 14 9 18 151 8 297 300 NOR2_X1 $T=55340 1000 0 0 $X=55225 $Y=885
X1909 13 9 34 291 8 297 300 NOR2_X1 $T=57810 1000 1 180 $X=57125 $Y=885
X1910 12 9 19 209 8 299 300 NOR2_X1 $T=58000 3800 0 180 $X=57315 $Y=2285
X1911 21 9 67 153 8 298 301 NOR2_X1 $T=57810 6600 1 0 $X=57695 $Y=5085
X1912 20 9 35 210 8 298 301 NOR2_X1 $T=58950 6600 0 180 $X=58265 $Y=5085
X1913 36 9 3 211 8 298 301 NOR2_X1 $T=59520 6600 0 180 $X=58835 $Y=5085
X1914 21 9 34 152 8 299 300 NOR2_X1 $T=59710 3800 1 0 $X=59595 $Y=2285
X1915 20 9 18 179 8 298 122 NOR2_X1 $T=60090 6600 0 0 $X=59975 $Y=6485
X1916 20 9 19 237 8 299 301 NOR2_X1 $T=60660 3800 0 0 $X=60545 $Y=3685
X1917 36 9 34 154 8 298 122 NOR2_X1 $T=60660 6600 0 0 $X=60545 $Y=6485
X1918 36 9 69 238 8 299 301 NOR2_X1 $T=61230 3800 0 0 $X=61115 $Y=3685
X1919 21 9 18 180 8 297 300 NOR2_X1 $T=61990 1000 0 0 $X=61875 $Y=885
X1920 36 9 18 280 8 298 301 NOR2_X1 $T=63510 6600 0 180 $X=62825 $Y=5085
X1921 36 9 19 157 8 298 301 NOR2_X1 $T=63510 6600 1 0 $X=63395 $Y=5085
X1922 20 9 34 214 8 298 122 NOR2_X1 $T=64460 6600 1 180 $X=63775 $Y=6485
X1923 180 9 155 239 8 297 300 NOR2_X1 $T=64840 1000 1 180 $X=64155 $Y=885
X1924 94 9 18 159 8 298 122 NOR2_X1 $T=65790 6600 0 0 $X=65675 $Y=6485
X1925 21 9 19 162 8 298 301 NOR2_X1 $T=68830 6600 1 0 $X=68715 $Y=5085
X1926 36 9 30 221 8 298 301 NOR2_X1 $T=70920 6600 1 0 $X=70805 $Y=5085
X1927 20 9 69 263 8 298 301 NOR2_X1 $T=71490 6600 1 0 $X=71375 $Y=5085
X1928 21 9 69 164 8 298 301 NOR2_X1 $T=74530 6600 0 180 $X=73845 $Y=5085
X1929 20 9 30 241 8 298 301 NOR2_X1 $T=75480 6600 1 0 $X=75365 $Y=5085
X1930 36 9 37 226 8 298 301 NOR2_X1 $T=76050 6600 1 0 $X=75935 $Y=5085
X1931 267 9 165 227 8 297 300 NOR2_X1 $T=78140 1000 0 0 $X=78025 $Y=885
X1932 228 9 169 175 8 298 301 NOR2_X1 $T=79090 6600 1 0 $X=78975 $Y=5085
X1933 21 9 30 174 8 299 300 NOR2_X1 $T=82320 3800 1 0 $X=82205 $Y=2285
X1934 20 9 37 244 8 299 301 NOR2_X1 $T=83460 3800 0 0 $X=83345 $Y=3685
X1935 36 9 4 245 8 299 301 NOR2_X1 $T=84030 3800 0 0 $X=83915 $Y=3685
X1936 99 9 73 230 8 298 122 NOR2_X1 $T=84220 6600 0 0 $X=84105 $Y=6485
X1937 8 215 281 240 9 299 301 XNOR2_X1 $T=65600 3800 0 0 $X=65485 $Y=3685
X1938 9 156 293 259 8 299 301 XOR2_X1 $T=63700 3800 1 180 $X=62445 $Y=3685
X1939 9 261 262 163 8 297 300 XOR2_X1 $T=70350 1000 0 0 $X=70235 $Y=885
X1940 9 264 223 262 8 297 300 XOR2_X1 $T=71490 1000 0 0 $X=71375 $Y=885
X1941 9 170 224 266 8 297 300 XOR2_X1 $T=74720 1000 0 0 $X=74605 $Y=885
X1942 9 229 225 242 8 299 300 XOR2_X1 $T=79850 3800 0 180 $X=78595 $Y=2285
X1943 214 8 280 156 9 298 122 NAND2_X1 $T=63890 6600 1 180 $X=63205 $Y=6485
X1944 180 8 155 213 9 297 300 NAND2_X1 $T=64270 1000 1 180 $X=63585 $Y=885
X1945 217 8 218 264 9 297 300 NAND2_X1 $T=66930 1000 0 0 $X=66815 $Y=885
X1946 216 8 158 218 9 299 300 NAND2_X1 $T=67500 3800 0 180 $X=66815 $Y=2285
X1947 267 8 165 173 9 297 300 NAND2_X1 $T=78140 1000 1 180 $X=77455 $Y=885
X1948 228 8 169 172 9 298 301 NAND2_X1 $T=79660 6600 1 0 $X=79545 $Y=5085
X1949 213 156 215 239 8 9 299 300 AOI21_X1 $T=63700 3800 1 0 $X=63585 $Y=2285
X1950 228 169 242 175 8 9 299 301 AOI21_X1 $T=79280 3800 0 0 $X=79165 $Y=3685
X1951 173 170 229 227 8 9 297 300 AOI21_X1 $T=79850 1000 0 0 $X=79735 $Y=885
X1952 283 172 106 175 8 9 298 301 AOI21_X1 $T=81370 6600 1 0 $X=81255 $Y=5085
X1953 172 173 243 171 8 9 299 301 AOI21_X1 $T=82510 3800 1 180 $X=81635 $Y=3685
X1957 100 123 182 231 9 8 284 299 300 FA_X1 $T=1000 3800 1 0 $X=885 $Y=2285
X1958 39 124 284 295 9 8 40 299 301 FA_X1 $T=1000 3800 0 0 $X=885 $Y=3685
X1959 231 111 74 57 9 8 183 298 122 FA_X1 $T=1000 6600 0 0 $X=885 $Y=6485
X1960 182 125 246 270 9 8 127 299 301 FA_X1 $T=4040 3800 0 0 $X=3925 $Y=3685
X1961 123 126 232 185 9 8 184 297 300 FA_X1 $T=4990 1000 0 0 $X=4875 $Y=885
X1962 124 127 183 58 9 8 41 298 301 FA_X1 $T=4990 6600 1 0 $X=4875 $Y=5085
X1963 42 247 77 184 9 8 75 298 122 FA_X1 $T=12020 6600 1 180 $X=8865 $Y=6485
X1964 295 128 78 186 9 8 247 297 300 FA_X1 $T=9170 1000 0 0 $X=9055 $Y=885
X1965 101 285 286 271 9 8 188 298 301 FA_X1 $T=12020 6600 1 0 $X=11905 $Y=5085
X1966 186 129 233 189 9 8 131 297 300 FA_X1 $T=12210 1000 0 0 $X=12095 $Y=885
X1967 79 1 80 62 9 8 272 298 122 FA_X1 $T=13350 6600 0 0 $X=13235 $Y=6485
X1968 102 131 188 272 9 8 187 298 301 FA_X1 $T=18100 6600 0 180 $X=14945 $Y=5085
X1969 128 130 249 190 9 8 248 297 300 FA_X1 $T=15250 1000 0 0 $X=15135 $Y=885
X1970 190 112 81 63 9 8 82 298 122 FA_X1 $T=16390 6600 0 0 $X=16275 $Y=6485
X1971 43 248 23 64 9 8 176 298 301 FA_X1 $T=18100 6600 1 0 $X=17985 $Y=5085
X1972 83 176 187 273 9 8 11 298 122 FA_X1 $T=19430 6600 0 0 $X=19315 $Y=6485
X1973 130 132 191 274 9 8 84 299 300 FA_X1 $T=19810 3800 1 0 $X=19695 $Y=2285
X1974 44 296 194 55 9 8 250 299 301 FA_X1 $T=22850 3800 0 0 $X=22735 $Y=3685
X1975 249 133 251 192 9 8 45 297 300 FA_X1 $T=23040 1000 0 0 $X=22925 $Y=885
X1976 273 134 250 65 9 8 46 298 122 FA_X1 $T=26270 6600 0 0 $X=26155 $Y=6485
X1977 296 135 287 195 9 8 193 297 300 FA_X1 $T=26650 1000 0 0 $X=26535 $Y=885
X1978 134 136 193 252 9 8 27 298 301 FA_X1 $T=27980 6600 1 0 $X=27865 $Y=5085
X1979 85 2 288 66 9 8 136 298 122 FA_X1 $T=29310 6600 0 0 $X=29195 $Y=6485
X1980 194 137 289 275 9 8 252 299 301 FA_X1 $T=30450 3800 0 0 $X=30335 $Y=3685
X1981 32 139 197 196 9 8 253 297 300 FA_X1 $T=38240 1000 1 180 $X=35085 $Y=885
X1982 86 138 177 70 9 8 141 298 122 FA_X1 $T=35770 6600 0 0 $X=35655 $Y=6485
X1983 276 140 198 199 9 8 144 299 301 FA_X1 $T=40330 3800 1 180 $X=37175 $Y=3685
X1984 87 113 110 276 9 8 201 298 122 FA_X1 $T=38810 6600 0 0 $X=38695 $Y=6485
X1985 88 141 253 254 9 8 203 299 301 FA_X1 $T=40330 3800 0 0 $X=40215 $Y=3685
X1986 103 143 200 202 9 8 254 297 300 FA_X1 $T=43560 1000 1 180 $X=40405 $Y=885
X1987 47 142 204 201 9 8 290 298 122 FA_X1 $T=41850 6600 0 0 $X=41735 $Y=6485
X1988 142 144 206 56 9 8 48 299 301 FA_X1 $T=43370 3800 0 0 $X=43255 $Y=3685
X1989 143 145 255 205 9 8 206 297 300 FA_X1 $T=43560 1000 0 0 $X=43445 $Y=885
X1990 204 146 89 107 9 8 150 298 122 FA_X1 $T=44890 6600 0 0 $X=44775 $Y=6485
X1991 104 147 207 278 9 8 146 298 301 FA_X1 $T=46980 6600 1 0 $X=46865 $Y=5085
X1992 50 148 290 203 9 8 49 298 122 FA_X1 $T=50970 6600 1 180 $X=47815 $Y=6485
X1993 91 149 208 277 9 8 90 299 300 FA_X1 $T=51160 3800 0 180 $X=48005 $Y=2285
X1994 148 150 178 279 9 8 51 298 122 FA_X1 $T=50970 6600 0 0 $X=50855 $Y=6485
X1995 149 234 235 236 9 8 256 297 300 FA_X1 $T=52300 1000 0 0 $X=52185 $Y=885
X1996 208 151 291 209 9 8 257 299 300 FA_X1 $T=54390 3800 1 0 $X=54275 $Y=2285
X1997 279 5 256 257 9 8 52 299 301 FA_X1 $T=57620 3800 1 180 $X=54465 $Y=3685
X1998 178 108 258 114 9 8 92 298 122 FA_X1 $T=57050 6600 0 0 $X=56935 $Y=6485
X1999 53 153 210 211 9 8 258 299 301 FA_X1 $T=60660 3800 1 180 $X=57505 $Y=3685
X2000 161 152 237 238 9 8 158 297 300 FA_X1 $T=58950 1000 0 0 $X=58835 $Y=885
X2001 260 160 95 115 9 8 220 298 122 FA_X1 $T=66360 6600 0 0 $X=66245 $Y=6485
X2002 282 162 263 221 9 8 261 299 301 FA_X1 $T=71300 3800 0 0 $X=71185 $Y=3685
X2003 265 6 260 282 9 8 165 298 122 FA_X1 $T=72820 6600 0 0 $X=72705 $Y=6485
X2004 166 164 241 226 9 8 167 299 301 FA_X1 $T=74340 3800 0 0 $X=74225 $Y=3685
X2005 97 166 109 71 9 8 268 298 122 FA_X1 $T=75860 6600 0 0 $X=75745 $Y=6485
X2006 54 268 269 72 9 8 169 298 122 FA_X1 $T=81940 6600 1 180 $X=78785 $Y=6485
X2007 105 174 244 245 9 8 269 297 300 FA_X1 $T=81750 1000 0 0 $X=81635 $Y=885
X2008 264 222 8 170 261 163 9 297 300 OAI22_X1 $T=72630 1000 0 0 $X=72515 $Y=885
X2009 280 9 292 293 8 93 298 122 NOR3_X1 $T=63320 6600 1 180 $X=62445 $Y=6485
X2010 170 9 227 171 8 181 299 301 NOR3_X1 $T=80990 3800 0 0 $X=80875 $Y=3685
X2011 281 9 223 224 225 96 8 299 300 NOR4_X1 $T=72630 3800 1 0 $X=72515 $Y=2285
X2012 181 9 243 230 22 98 8 298 122 NOR4_X1 $T=81940 6600 0 0 $X=81825 $Y=6485
X2013 73 7 175 8 9 171 298 301 OR3_X1 $T=84790 6600 0 180 $X=83725 $Y=5085
.ENDS
***************************************
.SUBCKT FloatingPointMultiplierSingle VSS VDD result[31] result[29] result[28] result[27] result[26] result[23] result[25] result[24] result[22] result[21] inputB[16] result[20] result[19] inputB[11] inputB[14] reset result[18] inputA[14]
+ inputA[13] inputA[8] inputA[10] inputA[11] inputA[12] inputA[9] inputA[6] result[17] result[16] result[15] result[14] result[13] result[12] en result[11] clk inputB[31] inputB[29] inputA[31] inputB[24]
+ inputB[30] inputA[25] inputA[26] inputA[27] inputA[24] inputA[28] inputA[16] inputB[13] inputB[10] inputB[9] inputB[8] inputA[7] inputB[5] inputB[3] inputA[0] inputA[3] inputA[2] inputA[1] result[30] result[6]
+ result[10] result[9] result[4] result[8] result[1] result[7] inputB[27] inputB[28] inputB[26] inputB[23] OF result[5] result[3] result[0] result[2] inputA[19] inputB[22] inputB[19] inputB[17] inputB[25]
+ inputA[17] inputB[21] inputA[30] inputA[20] inputA[23] inputB[20] inputA[29] inputA[22] inputA[18] inputB[6] inputB[15] inputA[21] inputA[15] inputB[18] inputB[12] inputA[4] inputB[4] inputA[5] inputB[7] inputB[1]
+ inputB[2] inputB[0] 901 902 903 904
** N=926 EP=106 IP=2416 FDC=23054
X0 76 5 14 24 786 25 35 inputA[13] inputA[14] inputA[10] inputA[8] inputA[12] inputA[11] inputA[9] inputA[6] 788 789 61 62 55
+ 58 63 69 67 65 reset clk VDD result[23] result[24] result[21] result[20] 44 result[17] 73 VSS result[13] en 78 result[30]
+ 22 result[25] 27 37 result[18] 160 46 40 59 result[14] result[11] result[10] result[31] 8 57 71 result[6] result[9] result[29] result[28]
+ result[27] result[26] result[22] result[19] result[16] result[15] result[12] 787 49 790 74 906 6 9 11 13 15 20 21 785
+ 26 28 31 36 43 50 42 70 80 60 917
+ ICV_6 $T=0 0 0 0 $X=0 $Y=79285
X1 inputB[31] 84 86 87 88 91 793 99 102 25 109 111 107 110 112 907 108 113 35 115
+ 116 117 114 795 118 125 130 128 131 133 141 143 798 797 148 74 76 VDD VSS 27
+ 71 73 OF 5 6 792 92 169 100 14 22 786 28 788 121 119 796 122 49 129
+ 137 146 result[1] 711 147 result[8] result[4] result[7] 85 40 80 result[2] 9 11 24 106 26 31 36 83
+ 120 61 126 50 59 58 62 60 136 138 63 65 150 152 151 104 96 98 101 reset
+ 127 135 139 140 142 144 145 790 149 710 90 13 93 15 21 789 43 123 124 132
+ 134 69 70 20 785 55 94 97 105 794 89 103 918 917
+ ICV_8 $T=0 0 0 0 $X=0 $Y=73640
X2 inputA[31] inputB[29] inputB[28] 159 35 84 inputB[30] inputB[26] inputB[27] inputB[25] 161 163 inputA[25] VSS inputB[24] 906 inputB[23] 90 792 67
+ 94 91 88 97 170 92 173 800 174 802 108 175 107 805 inputB[16] inputB[14] inputB[11] 795 189 123
+ 128 912 203 212 136 721 227 231 223 797 226 311 145 312 235 148 234 238 239 76
+ 236 247 252 815 816 819 160 VDD 169 99 96 102 105 799 187 120 124 193 125 214
+ 137 138 241 255 144 83 85 95 793 93 101 801 166 791 188 129 126 135 201 204
+ 210 224 232 818 812 149 179 168 178 192 908 result[0] result[5] result[3] 158 162 165 167 787 44
+ 42 150 151 152 254 156 89 103 104 177 106 109 127 130 133 218 140 142 143 229
+ 190 202 213 100 176 180 184 185 117 195 191 215 216 225 245 243 246 242 248 253
+ 249 803 804 182 796 118 122 198 208 221 147 237 250 86 710 87 98 794 119 132
+ 134 139 141 146 798 172 186 807 808 911 197 200 809 205 206 301 302 220 810 230
+ 171 196 181 183 806 194 199 211 207 222 217 219 228 811 233 813 240 244 814 251
+ 817 918 919
+ ICV_10 $T=0 0 0 0 $X=0 $Y=62485
X3 inputA[30] inputB[19] inputA[22] inputA[28] inputA[29] inputA[27] inputB[17] inputA[19] 262 inputA[26] 35 inputA[24] 84 170 821 inputA[23] 268 264 270 857
+ 282 176 283 299 488 308 307 233 733 331 VDD VSS 266 265 823 278 279 175 280 287
+ 288 290 286 271 323 284 328 326 356 319 209 314 160 167 417 273 804 352 359 806
+ 295 329 316 208 217 228 811 364 inputB[22] 315 78 267 732 486 296 827 324 269 259 158
+ 163 261 165 802 172 801 907 803 808 189 912 297 205 206 829 221 226 230 812 813
+ 239 237 240 242 245 250 330 272 824 294 317 322 276 281 368 444 313 361 318 320
+ 831 300 159 161 162 83 820 166 799 173 800 110 805 181 186 190 193 191 197 198
+ 809 212 213 828 215 721 222 830 229 235 249 327 246 815 252 816 254 253 325 819
+ 171 177 111 201 203 220 810 232 244 275 291 292 298 305 309 303 274 285 826 310
+ 263 731 277 289 825 293 389 304 321 822 814 306 919 920
+ ICV_11 $T=0 0 0 0 $X=0 $Y=56885
X4 inputB[21] inputB[20] 84 inputA[20] 261 35 259 822 340 342 334 346 732 835 349 179 441 363 838 842
+ 827 211 320 464 847 387 382 391 848 745 396 324 405 VDD VSS 262 276 272 265 271
+ 821 266 319 417 339 347 355 131 361 300 194 461 370 362 357 306 369 746 328 323
+ 359 264 416 267 336 420 280 329 183 824 825 294 366 199 356 297 843 373 376 829
+ 400 379 304 386 227 392 399 248 286 488 406 160 742 338 345 351 743 365 402 832
+ 168 112 747 263 335 337 275 358 435 911 364 200 202 299 207 210 302 308 307 309
+ 311 312 224 733 234 243 315 317 318 831 404 384 820 269 341 422 348 284 354 834
+ 290 840 844 378 380 828 401 846 388 377 316 385 330 83 344 350 281 353 114 837
+ 744 184 367 192 908 845 214 381 303 383 231 390 403 397 398 849 352 209 326 295
+ 731 274 283 823 113 285 293 195 305 310 327 325 429 187 839 371 393 395 296 270
+ 343 287 841 372 375 374 850 394 268 836 282 833 360 238 920 921
+ ICV_12 $T=0 0 0 0 $X=0 $Y=51285
X5 inputB[15] inputA[16] 84 inputA[17] 35 inputA[21] inputA[18] inputB[5] 343 755 423 425 422 426 427 354 428 432 424 757
+ 385 366 859 451 450 455 457 437 464 463 440 746 404 VDD VSS 412 477 417 340 434
+ 355 356 400 758 842 413 377 374 375 376 438 381 439 488 83 913 832 160 272 263
+ 414 852 834 855 347 856 348 835 836 837 436 99 399 420 336 362 845 301 380 452
+ 204 445 225 219 846 388 459 465 390 514 405 271 251 817 474 331 288 759 inputB[18] 116
+ 353 505 825 337 479 418 169 341 278 360 841 368 826 298 847 848 389 386 393 236
+ 460 394 850 247 421 853 858 442 466 472 335 264 415 756 338 379 351 433 370 46
+ 57 461 449 218 448 446 401 471 468 454 359 862 300 361 467 267 431 269 430 276
+ 352 854 358 8 121 37 839 371 372 373 443 447 830 456 387 745 395 313 357 818
+ 398 469 849 403 321 475 406 833 174 277 349 115 350 744 838 840 844 378 216 314
+ 397 742 851 342 453 383 458 402 473 419 861 470 743 363 843 462 747 860 921 922
+ ICV_13 $T=0 0 0 0 $X=0 $Y=45685
X6 inputB[6] inputA[15] inputB[3] 84 913 35 inputA[7] inputA[5] inputA[4] 851 inputB[4] 764 444 863 854 423 855 872 490 496
+ 866 265 506 869 VDD VSS 415 160 323 416 294 417 853 756 857 345 426 483 858 271
+ 188 489 185 448 359 377 336 379 500 511 326 401 862 461 512 440 515 469 472 471
+ 284 83 418 413 464 856 288 439 491 446 442 499 465 319 286 352 510 356 504 300
+ 860 420 507 475 362 369 357 385 364 759 914 493 320 466 480 412 495 449 765 346
+ 430 431 485 291 365 367 492 514 447 453 503 468 864 414 384 484 488 498 867 295
+ 361 868 370 399 316 328 755 478 419 421 428 156 178 433 482 436 57 859 443 451
+ 400 455 456 508 509 457 458 392 513 463 438 467 861 322 209 329 427 429 865 460
+ 497 501 502 474 481 432 758 494 396 487 435 923 922
+ ICV_14 $T=0 0 0 0 $X=0 $Y=40085
X7 inputB[10] inputB[9] inputB[13] inputB[12] inputB[7] 84 inputB[0] inputB[2] inputB[8] inputB[1] 520 438 523 182 870 35 480 493 inputA[1] 499
+ 464 inputA[0] 544 inputA[3] inputA[2] 554 557 559 502 562 503 563 573 514 581 VDD VSS 83 444 530
+ 412 764 265 336 271 417 413 479 286 771 273 348 488 425 532 369 326 487 536 357
+ 292 399 491 385 328 160 400 288 284 775 454 867 511 568 507 439 470 440 518 528
+ 519 517 909 477 525 524 481 420 915 871 37 484 486 196 356 329 370 362 461 437
+ 549 295 323 320 352 498 401 473 452 391 510 364 377 869 465 572 777 209 579 582
+ 765 561 478 534 540 567 569 576 577 791 384 379 863 852 529 117 807 490 543 546
+ 553 513 509 255 570 462 874 776 575 571 580 877 583 345 558 910 535 300 361 316
+ 773 556 774 564 508 566 515 876 778 359 495 496 866 770 415 279 864 319 344 339
+ 757 289 542 545 868 560 873 382 505 565 459 574 865 424 494 501 497 506 522 527
+ 482 916 533 914 537 548 875 516 769 538 500 521 526 485 492 541 772 550 555 512
+ 504 578 539 531 923 924
+ ICV_16 $T=0 0 0 0 $X=0 $Y=28885
X8 517 84 584 357 590 771 591 420 598 438 538 326 328 886 553 613 887 612 450 614
+ 562 284 620 874 577 507 640 580 642 892 VSS VDD 589 522 336 520 413 356 879 526
+ 423 530 872 882 533 417 599 600 286 399 558 323 544 401 320 773 549 555 440 559
+ 465 774 564 359 361 618 626 625 571 634 519 587 265 319 878 770 592 461 352 905
+ 329 271 178 316 180 602 370 400 46 514 510 616 511 560 615 617 888 488 621 209
+ 362 439 776 288 629 632 574 628 633 891 636 638 595 385 582 369 881 619 622 631
+ 890 635 639 518 516 300 916 535 489 608 772 910 445 876 641 585 596 543 777 880
+ 437 156 884 364 464 295 624 576 499 583 588 334 521 523 483 528 434 529 441 545
+ 607 548 610 775 563 565 223 377 627 573 572 778 769 527 554 550 557 556 561 889
+ 875 578 637 581 623 524 593 597 536 540 546 611 567 570 566 630 586 525 37 594
+ 532 883 601 603 605 885 609 873 568 575 579 877 347 606 924 925
+ ICV_17 $T=0 0 0 0 $X=0 $Y=19085
X9 894 589 649 652 319 660 882 539 599 514 465 464 679 685 499 636 891 635 705 700
+ 584 422 VSS VDD 271 438 329 286 336 265 594 361 915 316 357 400 420 488 377 288
+ 295 284 542 359 323 440 886 369 686 687 619 401 510 695 629 646 645 437 905 896
+ 300 854 909 779 370 664 669 413 670 188 8 399 672 356 611 507 511 328 689 690
+ 693 623 627 691 631 784 320 698 704 701 702 703 893 461 657 662 666 674 681 694
+ 783 870 643 590 895 656 593 653 663 596 531 595 537 600 884 541 606 885 781 612
+ 615 888 688 617 621 620 626 624 630 696 637 699 655 534 676 608 683 641 878 121
+ 352 417 667 385 362 898 209 364 439 675 326 610 622 569 625 644 587 591 871 592
+ 880 654 658 598 668 602 671 603 780 677 692 890 628 241 634 633 892 638 585 586
+ 588 156 607 605 609 613 887 616 640 642 614 618 648 650 528 673 678 782 889 632
+ 697 639 680 879 651 661 881 665 897 46 899 682 684 900 647 659 925 926
+ ICV_19 $T=0 0 0 0 $X=0 $Y=7885
X10 654 668 357 359 686 783 704 VSS VDD 323 597 361 300 356 329 499 320 507 510 702
+ 666 437 438 326 601 286 400 209 385 898 399 401 370 511 295 700 894 644 649 648
+ 651 659 665 883 899 680 679 681 684 685 683 698 663 687 645 647 464 420 413 657
+ 662 664 669 670 369 352 364 672 784 696 703 646 650 461 895 653 896 656 779 660
+ 661 897 667 671 676 673 781 682 782 690 691 465 693 695 697 705 701 893 652 655
+ 675 678 900 699 677 689 694 780 643 658 674 688 692 926
+ ICV_20 $T=0 0 0 0 $X=0 $Y=0
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
